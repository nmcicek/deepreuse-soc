  
module ArtixMMCM(
    input clk_in1_p,
    input clk_in1_n,
    output clk_out1,
    input reset,
    output locked
);

endmodule