module Queue_64( // @[:boom.system.TestHarness.MegaBoomConfig.fir@16911.2]
  input         clock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@16912.4]
  input         reset, // @[:boom.system.TestHarness.MegaBoomConfig.fir@16913.4]
  output        io_enq_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@16914.4]
  input         io_enq_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@16914.4]
  input  [15:0] io_enq_bits, // @[:boom.system.TestHarness.MegaBoomConfig.fir@16914.4]
  input         io_deq_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@16914.4]
  output        io_deq_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@16914.4]
  output [15:0] io_deq_bits // @[:boom.system.TestHarness.MegaBoomConfig.fir@16914.4]
);
  reg [15:0] _T_35 [0:15]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
  reg [31:0] _RAND_0;
  wire [15:0] _T_35__T_58_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
  wire [3:0] _T_35__T_58_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
  wire [15:0] _T_35__T_50_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
  wire [3:0] _T_35__T_50_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
  wire  _T_35__T_50_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
  wire  _T_35__T_50_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
  reg [3:0] value; // @[Counter.scala 26:33:boom.system.TestHarness.MegaBoomConfig.fir@16920.4]
  reg [31:0] _RAND_1;
  reg [3:0] value_1; // @[Counter.scala 26:33:boom.system.TestHarness.MegaBoomConfig.fir@16921.4]
  reg [31:0] _RAND_2;
  reg  _T_39; // @[Decoupled.scala 217:35:boom.system.TestHarness.MegaBoomConfig.fir@16922.4]
  reg [31:0] _RAND_3;
  wire  _T_40; // @[Decoupled.scala 219:41:boom.system.TestHarness.MegaBoomConfig.fir@16923.4]
  wire  _T_41; // @[Decoupled.scala 220:36:boom.system.TestHarness.MegaBoomConfig.fir@16924.4]
  wire  _T_42; // @[Decoupled.scala 220:33:boom.system.TestHarness.MegaBoomConfig.fir@16925.4]
  wire  _T_43; // @[Decoupled.scala 221:32:boom.system.TestHarness.MegaBoomConfig.fir@16926.4]
  wire  _T_44; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@16927.4]
  wire  _T_47; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@16931.4]
  wire [3:0] _T_52; // @[Counter.scala 35:22:boom.system.TestHarness.MegaBoomConfig.fir@16940.6]
  wire [3:0] _T_54; // @[Counter.scala 35:22:boom.system.TestHarness.MegaBoomConfig.fir@16946.6]
  wire  _T_55; // @[Decoupled.scala 232:16:boom.system.TestHarness.MegaBoomConfig.fir@16949.4]
  assign _T_35__T_58_addr = value_1;
  assign _T_35__T_58_data = _T_35[_T_35__T_58_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
  assign _T_35__T_50_data = io_enq_bits;
  assign _T_35__T_50_addr = value;
  assign _T_35__T_50_mask = 1'h1;
  assign _T_35__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_40 = value == value_1; // @[Decoupled.scala 219:41:boom.system.TestHarness.MegaBoomConfig.fir@16923.4]
  assign _T_41 = _T_39 == 1'h0; // @[Decoupled.scala 220:36:boom.system.TestHarness.MegaBoomConfig.fir@16924.4]
  assign _T_42 = _T_40 & _T_41; // @[Decoupled.scala 220:33:boom.system.TestHarness.MegaBoomConfig.fir@16925.4]
  assign _T_43 = _T_40 & _T_39; // @[Decoupled.scala 221:32:boom.system.TestHarness.MegaBoomConfig.fir@16926.4]
  assign _T_44 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@16927.4]
  assign _T_47 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@16931.4]
  assign _T_52 = value + 4'h1; // @[Counter.scala 35:22:boom.system.TestHarness.MegaBoomConfig.fir@16940.6]
  assign _T_54 = value_1 + 4'h1; // @[Counter.scala 35:22:boom.system.TestHarness.MegaBoomConfig.fir@16946.6]
  assign _T_55 = _T_44 != _T_47; // @[Decoupled.scala 232:16:boom.system.TestHarness.MegaBoomConfig.fir@16949.4]
  assign io_enq_ready = _T_43 == 1'h0; // @[Decoupled.scala 237:16:boom.system.TestHarness.MegaBoomConfig.fir@16956.4]
  assign io_deq_valid = _T_42 == 1'h0; // @[Decoupled.scala 236:16:boom.system.TestHarness.MegaBoomConfig.fir@16954.4]
  assign io_deq_bits = _T_35__T_58_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@16958.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    _T_35[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_39 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35__T_50_en & _T_35__T_50_mask) begin
      _T_35[_T_35__T_50_addr] <= _T_35__T_50_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@16919.4]
    end
    if (reset) begin
      value <= 4'h0;
    end else begin
      if (_T_44) begin
        value <= _T_52;
      end
    end
    if (reset) begin
      value_1 <= 4'h0;
    end else begin
      if (_T_47) begin
        value_1 <= _T_54;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_55) begin
        _T_39 <= _T_44;
      end
    end
  end
endmodule
module AXI4UserYanker_2( // @[:boom.system.TestHarness.MegaBoomConfig.fir@18671.2]
  input         clock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18672.4]
  input         reset, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18673.4]
  output        auto_in_aw_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_in_aw_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [3:0]  auto_in_aw_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [31:0] auto_in_aw_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_in_aw_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [15:0] auto_in_aw_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_in_w_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_in_w_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [63:0] auto_in_w_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [7:0]  auto_in_w_bits_strb, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_in_w_bits_last, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_in_b_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_in_b_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [3:0]  auto_in_b_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [1:0]  auto_in_b_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [15:0] auto_in_b_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_in_ar_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_in_ar_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [3:0]  auto_in_ar_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [31:0] auto_in_ar_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_in_ar_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [15:0] auto_in_ar_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_in_r_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_in_r_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [3:0]  auto_in_r_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [63:0] auto_in_r_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [1:0]  auto_in_r_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [15:0] auto_in_r_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_in_r_bits_last, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_out_aw_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_out_aw_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [3:0]  auto_out_aw_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [31:0] auto_out_aw_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [7:0]  auto_out_aw_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [2:0]  auto_out_aw_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_out_aw_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_out_w_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_out_w_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [63:0] auto_out_w_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [7:0]  auto_out_w_bits_strb, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_out_w_bits_last, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_out_b_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_out_b_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [3:0]  auto_out_b_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_out_ar_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_out_ar_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [3:0]  auto_out_ar_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [31:0] auto_out_ar_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [7:0]  auto_out_ar_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [2:0]  auto_out_ar_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_out_ar_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  output        auto_out_r_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_out_r_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [3:0]  auto_out_r_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [63:0] auto_out_r_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
  input         auto_out_r_bits_last // @[:boom.system.TestHarness.MegaBoomConfig.fir@18674.4]
);
  wire  Queue_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
  wire  Queue_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
  wire  Queue_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
  wire  Queue_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
  wire [15:0] Queue_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
  wire  Queue_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
  wire  Queue_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
  wire [15:0] Queue_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
  wire  Queue_1_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
  wire  Queue_1_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
  wire  Queue_1_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
  wire  Queue_1_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
  wire [15:0] Queue_1_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
  wire  Queue_1_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
  wire  Queue_1_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
  wire [15:0] Queue_1_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
  wire  Queue_2_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
  wire  Queue_2_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
  wire  Queue_2_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
  wire  Queue_2_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
  wire [15:0] Queue_2_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
  wire  Queue_2_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
  wire  Queue_2_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
  wire [15:0] Queue_2_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
  wire  Queue_3_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
  wire  Queue_3_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
  wire  Queue_3_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
  wire  Queue_3_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
  wire [15:0] Queue_3_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
  wire  Queue_3_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
  wire  Queue_3_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
  wire [15:0] Queue_3_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
  wire  Queue_4_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
  wire  Queue_4_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
  wire  Queue_4_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
  wire  Queue_4_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
  wire [15:0] Queue_4_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
  wire  Queue_4_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
  wire  Queue_4_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
  wire [15:0] Queue_4_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
  wire  Queue_5_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
  wire  Queue_5_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
  wire  Queue_5_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
  wire  Queue_5_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
  wire [15:0] Queue_5_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
  wire  Queue_5_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
  wire  Queue_5_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
  wire [15:0] Queue_5_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
  wire  Queue_6_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
  wire  Queue_6_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
  wire  Queue_6_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
  wire  Queue_6_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
  wire [15:0] Queue_6_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
  wire  Queue_6_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
  wire  Queue_6_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
  wire [15:0] Queue_6_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
  wire  Queue_7_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
  wire  Queue_7_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
  wire  Queue_7_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
  wire  Queue_7_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
  wire [15:0] Queue_7_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
  wire  Queue_7_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
  wire  Queue_7_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
  wire [15:0] Queue_7_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
  wire  Queue_8_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
  wire  Queue_8_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
  wire  Queue_8_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
  wire  Queue_8_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
  wire [15:0] Queue_8_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
  wire  Queue_8_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
  wire  Queue_8_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
  wire [15:0] Queue_8_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
  wire  Queue_9_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
  wire  Queue_9_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
  wire  Queue_9_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
  wire  Queue_9_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
  wire [15:0] Queue_9_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
  wire  Queue_9_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
  wire  Queue_9_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
  wire [15:0] Queue_9_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
  wire  Queue_10_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
  wire  Queue_10_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
  wire  Queue_10_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
  wire  Queue_10_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
  wire [15:0] Queue_10_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
  wire  Queue_10_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
  wire  Queue_10_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
  wire [15:0] Queue_10_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
  wire  Queue_11_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
  wire  Queue_11_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
  wire  Queue_11_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
  wire  Queue_11_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
  wire [15:0] Queue_11_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
  wire  Queue_11_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
  wire  Queue_11_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
  wire [15:0] Queue_11_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
  wire  Queue_12_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
  wire  Queue_12_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
  wire  Queue_12_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
  wire  Queue_12_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
  wire [15:0] Queue_12_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
  wire  Queue_12_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
  wire  Queue_12_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
  wire [15:0] Queue_12_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
  wire  Queue_13_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
  wire  Queue_13_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
  wire  Queue_13_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
  wire  Queue_13_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
  wire [15:0] Queue_13_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
  wire  Queue_13_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
  wire  Queue_13_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
  wire [15:0] Queue_13_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
  wire  Queue_14_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
  wire  Queue_14_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
  wire  Queue_14_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
  wire  Queue_14_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
  wire [15:0] Queue_14_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
  wire  Queue_14_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
  wire  Queue_14_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
  wire [15:0] Queue_14_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
  wire  Queue_15_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
  wire  Queue_15_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
  wire  Queue_15_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
  wire  Queue_15_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
  wire [15:0] Queue_15_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
  wire  Queue_15_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
  wire  Queue_15_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
  wire [15:0] Queue_15_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
  wire  Queue_16_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
  wire  Queue_16_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
  wire  Queue_16_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
  wire  Queue_16_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
  wire [15:0] Queue_16_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
  wire  Queue_16_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
  wire  Queue_16_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
  wire [15:0] Queue_16_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
  wire  Queue_17_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
  wire  Queue_17_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
  wire  Queue_17_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
  wire  Queue_17_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
  wire [15:0] Queue_17_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
  wire  Queue_17_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
  wire  Queue_17_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
  wire [15:0] Queue_17_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
  wire  Queue_18_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
  wire  Queue_18_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
  wire  Queue_18_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
  wire  Queue_18_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
  wire [15:0] Queue_18_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
  wire  Queue_18_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
  wire  Queue_18_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
  wire [15:0] Queue_18_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
  wire  Queue_19_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
  wire  Queue_19_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
  wire  Queue_19_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
  wire  Queue_19_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
  wire [15:0] Queue_19_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
  wire  Queue_19_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
  wire  Queue_19_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
  wire [15:0] Queue_19_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
  wire  Queue_20_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
  wire  Queue_20_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
  wire  Queue_20_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
  wire  Queue_20_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
  wire [15:0] Queue_20_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
  wire  Queue_20_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
  wire  Queue_20_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
  wire [15:0] Queue_20_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
  wire  Queue_21_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
  wire  Queue_21_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
  wire  Queue_21_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
  wire  Queue_21_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
  wire [15:0] Queue_21_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
  wire  Queue_21_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
  wire  Queue_21_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
  wire [15:0] Queue_21_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
  wire  Queue_22_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
  wire  Queue_22_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
  wire  Queue_22_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
  wire  Queue_22_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
  wire [15:0] Queue_22_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
  wire  Queue_22_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
  wire  Queue_22_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
  wire [15:0] Queue_22_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
  wire  Queue_23_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
  wire  Queue_23_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
  wire  Queue_23_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
  wire  Queue_23_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
  wire [15:0] Queue_23_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
  wire  Queue_23_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
  wire  Queue_23_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
  wire [15:0] Queue_23_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
  wire  Queue_24_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
  wire  Queue_24_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
  wire  Queue_24_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
  wire  Queue_24_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
  wire [15:0] Queue_24_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
  wire  Queue_24_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
  wire  Queue_24_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
  wire [15:0] Queue_24_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
  wire  Queue_25_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
  wire  Queue_25_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
  wire  Queue_25_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
  wire  Queue_25_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
  wire [15:0] Queue_25_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
  wire  Queue_25_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
  wire  Queue_25_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
  wire [15:0] Queue_25_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
  wire  Queue_26_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
  wire  Queue_26_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
  wire  Queue_26_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
  wire  Queue_26_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
  wire [15:0] Queue_26_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
  wire  Queue_26_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
  wire  Queue_26_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
  wire [15:0] Queue_26_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
  wire  Queue_27_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
  wire  Queue_27_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
  wire  Queue_27_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
  wire  Queue_27_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
  wire [15:0] Queue_27_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
  wire  Queue_27_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
  wire  Queue_27_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
  wire [15:0] Queue_27_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
  wire  Queue_28_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
  wire  Queue_28_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
  wire  Queue_28_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
  wire  Queue_28_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
  wire [15:0] Queue_28_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
  wire  Queue_28_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
  wire  Queue_28_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
  wire [15:0] Queue_28_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
  wire  Queue_29_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
  wire  Queue_29_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
  wire  Queue_29_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
  wire  Queue_29_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
  wire [15:0] Queue_29_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
  wire  Queue_29_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
  wire  Queue_29_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
  wire [15:0] Queue_29_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
  wire  Queue_30_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
  wire  Queue_30_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
  wire  Queue_30_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
  wire  Queue_30_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
  wire [15:0] Queue_30_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
  wire  Queue_30_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
  wire  Queue_30_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
  wire [15:0] Queue_30_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
  wire  Queue_31_clock; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
  wire  Queue_31_reset; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
  wire  Queue_31_io_enq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
  wire  Queue_31_io_enq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
  wire [15:0] Queue_31_io_enq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
  wire  Queue_31_io_deq_ready; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
  wire  Queue_31_io_deq_valid; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
  wire [15:0] Queue_31_io_deq_bits; // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
  wire  _T_224_0; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18815.4]
  wire  _T_224_1; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18816.4]
  wire  _GEN_1; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_2; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18817.4]
  wire  _GEN_2; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_3; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18818.4]
  wire  _GEN_3; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_4; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18819.4]
  wire  _GEN_4; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_5; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18820.4]
  wire  _GEN_5; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_6; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18821.4]
  wire  _GEN_6; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_7; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18822.4]
  wire  _GEN_7; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_8; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18823.4]
  wire  _GEN_8; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_9; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18824.4]
  wire  _GEN_9; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_10; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18825.4]
  wire  _GEN_10; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_11; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18826.4]
  wire  _GEN_11; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_12; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18827.4]
  wire  _GEN_12; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_13; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18828.4]
  wire  _GEN_13; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_14; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18829.4]
  wire  _GEN_14; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_224_15; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18830.4]
  wire  _GEN_15; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  wire  _T_292; // @[UserYanker.scala 54:15:boom.system.TestHarness.MegaBoomConfig.fir@18872.4]
  wire  _T_249_0; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18838.4]
  wire  _T_249_1; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18839.4]
  wire  _GEN_17; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_2; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18840.4]
  wire  _GEN_18; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_3; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18841.4]
  wire  _GEN_19; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_4; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18842.4]
  wire  _GEN_20; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_5; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18843.4]
  wire  _GEN_21; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_6; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18844.4]
  wire  _GEN_22; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_7; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18845.4]
  wire  _GEN_23; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_8; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18846.4]
  wire  _GEN_24; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_9; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18847.4]
  wire  _GEN_25; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_10; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18848.4]
  wire  _GEN_26; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_11; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18849.4]
  wire  _GEN_27; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_12; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18850.4]
  wire  _GEN_28; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_13; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18851.4]
  wire  _GEN_29; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_14; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18852.4]
  wire  _GEN_30; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_249_15; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18853.4]
  wire  _GEN_31; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_293; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  wire  _T_295; // @[UserYanker.scala 54:14:boom.system.TestHarness.MegaBoomConfig.fir@18875.4]
  wire  _T_296; // @[UserYanker.scala 54:14:boom.system.TestHarness.MegaBoomConfig.fir@18876.4]
  wire [15:0] _T_272_0; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18856.4]
  wire [15:0] _T_272_1; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18857.4]
  wire [15:0] _GEN_33; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_2; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18858.4]
  wire [15:0] _GEN_34; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_3; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18859.4]
  wire [15:0] _GEN_35; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_4; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18860.4]
  wire [15:0] _GEN_36; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_5; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18861.4]
  wire [15:0] _GEN_37; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_6; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18862.4]
  wire [15:0] _GEN_38; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_7; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18863.4]
  wire [15:0] _GEN_39; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_8; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18864.4]
  wire [15:0] _GEN_40; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_9; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18865.4]
  wire [15:0] _GEN_41; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_10; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18866.4]
  wire [15:0] _GEN_42; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_11; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18867.4]
  wire [15:0] _GEN_43; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_12; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18868.4]
  wire [15:0] _GEN_44; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_13; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18869.4]
  wire [15:0] _GEN_45; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_14; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18870.4]
  wire [15:0] _GEN_46; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  wire [15:0] _T_272_15; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18871.4]
  wire [15:0] _T_298; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@18884.4]
  wire  _T_300; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18886.4]
  wire  _T_301; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18887.4]
  wire  _T_302; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18888.4]
  wire  _T_303; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18889.4]
  wire  _T_304; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18890.4]
  wire  _T_305; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18891.4]
  wire  _T_306; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18892.4]
  wire  _T_307; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18893.4]
  wire  _T_308; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18894.4]
  wire  _T_309; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18895.4]
  wire  _T_310; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18896.4]
  wire  _T_311; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18897.4]
  wire  _T_312; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18898.4]
  wire  _T_313; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18899.4]
  wire  _T_314; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18900.4]
  wire  _T_315; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18901.4]
  wire [15:0] _T_317; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@18903.4]
  wire  _T_319; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18905.4]
  wire  _T_320; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18906.4]
  wire  _T_321; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18907.4]
  wire  _T_322; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18908.4]
  wire  _T_323; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18909.4]
  wire  _T_324; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18910.4]
  wire  _T_325; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18911.4]
  wire  _T_326; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18912.4]
  wire  _T_327; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18913.4]
  wire  _T_328; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18914.4]
  wire  _T_329; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18915.4]
  wire  _T_330; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18916.4]
  wire  _T_331; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18917.4]
  wire  _T_332; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18918.4]
  wire  _T_333; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18919.4]
  wire  _T_334; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18920.4]
  wire  _T_335; // @[UserYanker.scala 61:37:boom.system.TestHarness.MegaBoomConfig.fir@18921.4]
  wire  _T_336; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18922.4]
  wire  _T_338; // @[UserYanker.scala 62:37:boom.system.TestHarness.MegaBoomConfig.fir@18925.4]
  wire  _T_341; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18930.4]
  wire  _T_346; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18938.4]
  wire  _T_351; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18946.4]
  wire  _T_356; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18954.4]
  wire  _T_361; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18962.4]
  wire  _T_366; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18970.4]
  wire  _T_371; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18978.4]
  wire  _T_376; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18986.4]
  wire  _T_381; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18994.4]
  wire  _T_386; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19002.4]
  wire  _T_391; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19010.4]
  wire  _T_396; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19018.4]
  wire  _T_401; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19026.4]
  wire  _T_406; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19034.4]
  wire  _T_411; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19042.4]
  wire  _T_418_0; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19051.4]
  wire  _T_418_1; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19052.4]
  wire  _GEN_49; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_2; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19053.4]
  wire  _GEN_50; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_3; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19054.4]
  wire  _GEN_51; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_4; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19055.4]
  wire  _GEN_52; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_5; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19056.4]
  wire  _GEN_53; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_6; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19057.4]
  wire  _GEN_54; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_7; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19058.4]
  wire  _GEN_55; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_8; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19059.4]
  wire  _GEN_56; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_9; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19060.4]
  wire  _GEN_57; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_10; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19061.4]
  wire  _GEN_58; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_11; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19062.4]
  wire  _GEN_59; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_12; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19063.4]
  wire  _GEN_60; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_13; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19064.4]
  wire  _GEN_61; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_14; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19065.4]
  wire  _GEN_62; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_418_15; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19066.4]
  wire  _GEN_63; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  wire  _T_486; // @[UserYanker.scala 75:15:boom.system.TestHarness.MegaBoomConfig.fir@19108.4]
  wire  _T_443_0; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19074.4]
  wire  _T_443_1; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19075.4]
  wire  _GEN_65; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_2; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19076.4]
  wire  _GEN_66; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_3; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19077.4]
  wire  _GEN_67; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_4; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19078.4]
  wire  _GEN_68; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_5; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19079.4]
  wire  _GEN_69; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_6; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19080.4]
  wire  _GEN_70; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_7; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19081.4]
  wire  _GEN_71; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_8; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19082.4]
  wire  _GEN_72; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_9; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19083.4]
  wire  _GEN_73; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_10; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19084.4]
  wire  _GEN_74; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_11; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19085.4]
  wire  _GEN_75; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_12; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19086.4]
  wire  _GEN_76; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_13; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19087.4]
  wire  _GEN_77; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_14; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19088.4]
  wire  _GEN_78; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_443_15; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19089.4]
  wire  _GEN_79; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_487; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  wire  _T_489; // @[UserYanker.scala 75:14:boom.system.TestHarness.MegaBoomConfig.fir@19111.4]
  wire  _T_490; // @[UserYanker.scala 75:14:boom.system.TestHarness.MegaBoomConfig.fir@19112.4]
  wire [15:0] _T_466_0; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19092.4]
  wire [15:0] _T_466_1; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19093.4]
  wire [15:0] _GEN_81; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_2; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19094.4]
  wire [15:0] _GEN_82; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_3; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19095.4]
  wire [15:0] _GEN_83; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_4; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19096.4]
  wire [15:0] _GEN_84; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_5; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19097.4]
  wire [15:0] _GEN_85; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_6; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19098.4]
  wire [15:0] _GEN_86; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_7; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19099.4]
  wire [15:0] _GEN_87; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_8; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19100.4]
  wire [15:0] _GEN_88; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_9; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19101.4]
  wire [15:0] _GEN_89; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_10; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19102.4]
  wire [15:0] _GEN_90; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_11; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19103.4]
  wire [15:0] _GEN_91; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_12; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19104.4]
  wire [15:0] _GEN_92; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_13; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19105.4]
  wire [15:0] _GEN_93; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_14; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19106.4]
  wire [15:0] _GEN_94; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  wire [15:0] _T_466_15; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19107.4]
  wire [15:0] _T_492; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@19120.4]
  wire  _T_494; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19122.4]
  wire  _T_495; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19123.4]
  wire  _T_496; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19124.4]
  wire  _T_497; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19125.4]
  wire  _T_498; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19126.4]
  wire  _T_499; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19127.4]
  wire  _T_500; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19128.4]
  wire  _T_501; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19129.4]
  wire  _T_502; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19130.4]
  wire  _T_503; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19131.4]
  wire  _T_504; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19132.4]
  wire  _T_505; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19133.4]
  wire  _T_506; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19134.4]
  wire  _T_507; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19135.4]
  wire  _T_508; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19136.4]
  wire  _T_509; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19137.4]
  wire [15:0] _T_511; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@19139.4]
  wire  _T_513; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19141.4]
  wire  _T_514; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19142.4]
  wire  _T_515; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19143.4]
  wire  _T_516; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19144.4]
  wire  _T_517; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19145.4]
  wire  _T_518; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19146.4]
  wire  _T_519; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19147.4]
  wire  _T_520; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19148.4]
  wire  _T_521; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19149.4]
  wire  _T_522; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19150.4]
  wire  _T_523; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19151.4]
  wire  _T_524; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19152.4]
  wire  _T_525; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19153.4]
  wire  _T_526; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19154.4]
  wire  _T_527; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19155.4]
  wire  _T_528; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19156.4]
  wire  _T_529; // @[UserYanker.scala 82:37:boom.system.TestHarness.MegaBoomConfig.fir@19157.4]
  wire  _T_531; // @[UserYanker.scala 83:37:boom.system.TestHarness.MegaBoomConfig.fir@19160.4]
  Queue_64 Queue ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18685.4]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  Queue_64 Queue_1 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18689.4]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  Queue_64 Queue_2 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18693.4]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  Queue_64 Queue_3 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18697.4]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  Queue_64 Queue_4 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18701.4]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits(Queue_4_io_enq_bits),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits(Queue_4_io_deq_bits)
  );
  Queue_64 Queue_5 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18705.4]
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits(Queue_5_io_enq_bits),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits(Queue_5_io_deq_bits)
  );
  Queue_64 Queue_6 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18709.4]
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits(Queue_6_io_enq_bits),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits(Queue_6_io_deq_bits)
  );
  Queue_64 Queue_7 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18713.4]
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits(Queue_7_io_enq_bits),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits(Queue_7_io_deq_bits)
  );
  Queue_64 Queue_8 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18717.4]
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits(Queue_8_io_enq_bits),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits(Queue_8_io_deq_bits)
  );
  Queue_64 Queue_9 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18721.4]
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits(Queue_9_io_enq_bits),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits(Queue_9_io_deq_bits)
  );
  Queue_64 Queue_10 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18725.4]
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits(Queue_10_io_enq_bits),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits(Queue_10_io_deq_bits)
  );
  Queue_64 Queue_11 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18729.4]
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits(Queue_11_io_enq_bits),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits(Queue_11_io_deq_bits)
  );
  Queue_64 Queue_12 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18733.4]
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits(Queue_12_io_enq_bits),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits(Queue_12_io_deq_bits)
  );
  Queue_64 Queue_13 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18737.4]
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits(Queue_13_io_enq_bits),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits(Queue_13_io_deq_bits)
  );
  Queue_64 Queue_14 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18741.4]
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits(Queue_14_io_enq_bits),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits(Queue_14_io_deq_bits)
  );
  Queue_64 Queue_15 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18745.4]
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits(Queue_15_io_enq_bits),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits(Queue_15_io_deq_bits)
  );
  Queue_64 Queue_16 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18749.4]
    .clock(Queue_16_clock),
    .reset(Queue_16_reset),
    .io_enq_ready(Queue_16_io_enq_ready),
    .io_enq_valid(Queue_16_io_enq_valid),
    .io_enq_bits(Queue_16_io_enq_bits),
    .io_deq_ready(Queue_16_io_deq_ready),
    .io_deq_valid(Queue_16_io_deq_valid),
    .io_deq_bits(Queue_16_io_deq_bits)
  );
  Queue_64 Queue_17 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18753.4]
    .clock(Queue_17_clock),
    .reset(Queue_17_reset),
    .io_enq_ready(Queue_17_io_enq_ready),
    .io_enq_valid(Queue_17_io_enq_valid),
    .io_enq_bits(Queue_17_io_enq_bits),
    .io_deq_ready(Queue_17_io_deq_ready),
    .io_deq_valid(Queue_17_io_deq_valid),
    .io_deq_bits(Queue_17_io_deq_bits)
  );
  Queue_64 Queue_18 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18757.4]
    .clock(Queue_18_clock),
    .reset(Queue_18_reset),
    .io_enq_ready(Queue_18_io_enq_ready),
    .io_enq_valid(Queue_18_io_enq_valid),
    .io_enq_bits(Queue_18_io_enq_bits),
    .io_deq_ready(Queue_18_io_deq_ready),
    .io_deq_valid(Queue_18_io_deq_valid),
    .io_deq_bits(Queue_18_io_deq_bits)
  );
  Queue_64 Queue_19 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18761.4]
    .clock(Queue_19_clock),
    .reset(Queue_19_reset),
    .io_enq_ready(Queue_19_io_enq_ready),
    .io_enq_valid(Queue_19_io_enq_valid),
    .io_enq_bits(Queue_19_io_enq_bits),
    .io_deq_ready(Queue_19_io_deq_ready),
    .io_deq_valid(Queue_19_io_deq_valid),
    .io_deq_bits(Queue_19_io_deq_bits)
  );
  Queue_64 Queue_20 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18765.4]
    .clock(Queue_20_clock),
    .reset(Queue_20_reset),
    .io_enq_ready(Queue_20_io_enq_ready),
    .io_enq_valid(Queue_20_io_enq_valid),
    .io_enq_bits(Queue_20_io_enq_bits),
    .io_deq_ready(Queue_20_io_deq_ready),
    .io_deq_valid(Queue_20_io_deq_valid),
    .io_deq_bits(Queue_20_io_deq_bits)
  );
  Queue_64 Queue_21 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18769.4]
    .clock(Queue_21_clock),
    .reset(Queue_21_reset),
    .io_enq_ready(Queue_21_io_enq_ready),
    .io_enq_valid(Queue_21_io_enq_valid),
    .io_enq_bits(Queue_21_io_enq_bits),
    .io_deq_ready(Queue_21_io_deq_ready),
    .io_deq_valid(Queue_21_io_deq_valid),
    .io_deq_bits(Queue_21_io_deq_bits)
  );
  Queue_64 Queue_22 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18773.4]
    .clock(Queue_22_clock),
    .reset(Queue_22_reset),
    .io_enq_ready(Queue_22_io_enq_ready),
    .io_enq_valid(Queue_22_io_enq_valid),
    .io_enq_bits(Queue_22_io_enq_bits),
    .io_deq_ready(Queue_22_io_deq_ready),
    .io_deq_valid(Queue_22_io_deq_valid),
    .io_deq_bits(Queue_22_io_deq_bits)
  );
  Queue_64 Queue_23 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18777.4]
    .clock(Queue_23_clock),
    .reset(Queue_23_reset),
    .io_enq_ready(Queue_23_io_enq_ready),
    .io_enq_valid(Queue_23_io_enq_valid),
    .io_enq_bits(Queue_23_io_enq_bits),
    .io_deq_ready(Queue_23_io_deq_ready),
    .io_deq_valid(Queue_23_io_deq_valid),
    .io_deq_bits(Queue_23_io_deq_bits)
  );
  Queue_64 Queue_24 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18781.4]
    .clock(Queue_24_clock),
    .reset(Queue_24_reset),
    .io_enq_ready(Queue_24_io_enq_ready),
    .io_enq_valid(Queue_24_io_enq_valid),
    .io_enq_bits(Queue_24_io_enq_bits),
    .io_deq_ready(Queue_24_io_deq_ready),
    .io_deq_valid(Queue_24_io_deq_valid),
    .io_deq_bits(Queue_24_io_deq_bits)
  );
  Queue_64 Queue_25 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18785.4]
    .clock(Queue_25_clock),
    .reset(Queue_25_reset),
    .io_enq_ready(Queue_25_io_enq_ready),
    .io_enq_valid(Queue_25_io_enq_valid),
    .io_enq_bits(Queue_25_io_enq_bits),
    .io_deq_ready(Queue_25_io_deq_ready),
    .io_deq_valid(Queue_25_io_deq_valid),
    .io_deq_bits(Queue_25_io_deq_bits)
  );
  Queue_64 Queue_26 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18789.4]
    .clock(Queue_26_clock),
    .reset(Queue_26_reset),
    .io_enq_ready(Queue_26_io_enq_ready),
    .io_enq_valid(Queue_26_io_enq_valid),
    .io_enq_bits(Queue_26_io_enq_bits),
    .io_deq_ready(Queue_26_io_deq_ready),
    .io_deq_valid(Queue_26_io_deq_valid),
    .io_deq_bits(Queue_26_io_deq_bits)
  );
  Queue_64 Queue_27 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18793.4]
    .clock(Queue_27_clock),
    .reset(Queue_27_reset),
    .io_enq_ready(Queue_27_io_enq_ready),
    .io_enq_valid(Queue_27_io_enq_valid),
    .io_enq_bits(Queue_27_io_enq_bits),
    .io_deq_ready(Queue_27_io_deq_ready),
    .io_deq_valid(Queue_27_io_deq_valid),
    .io_deq_bits(Queue_27_io_deq_bits)
  );
  Queue_64 Queue_28 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18797.4]
    .clock(Queue_28_clock),
    .reset(Queue_28_reset),
    .io_enq_ready(Queue_28_io_enq_ready),
    .io_enq_valid(Queue_28_io_enq_valid),
    .io_enq_bits(Queue_28_io_enq_bits),
    .io_deq_ready(Queue_28_io_deq_ready),
    .io_deq_valid(Queue_28_io_deq_valid),
    .io_deq_bits(Queue_28_io_deq_bits)
  );
  Queue_64 Queue_29 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18801.4]
    .clock(Queue_29_clock),
    .reset(Queue_29_reset),
    .io_enq_ready(Queue_29_io_enq_ready),
    .io_enq_valid(Queue_29_io_enq_valid),
    .io_enq_bits(Queue_29_io_enq_bits),
    .io_deq_ready(Queue_29_io_deq_ready),
    .io_deq_valid(Queue_29_io_deq_valid),
    .io_deq_bits(Queue_29_io_deq_bits)
  );
  Queue_64 Queue_30 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18805.4]
    .clock(Queue_30_clock),
    .reset(Queue_30_reset),
    .io_enq_ready(Queue_30_io_enq_ready),
    .io_enq_valid(Queue_30_io_enq_valid),
    .io_enq_bits(Queue_30_io_enq_bits),
    .io_deq_ready(Queue_30_io_deq_ready),
    .io_deq_valid(Queue_30_io_deq_valid),
    .io_deq_bits(Queue_30_io_deq_bits)
  );
  Queue_64 Queue_31 ( // @[UserYanker.scala 38:17:boom.system.TestHarness.MegaBoomConfig.fir@18809.4]
    .clock(Queue_31_clock),
    .reset(Queue_31_reset),
    .io_enq_ready(Queue_31_io_enq_ready),
    .io_enq_valid(Queue_31_io_enq_valid),
    .io_enq_bits(Queue_31_io_enq_bits),
    .io_deq_ready(Queue_31_io_deq_ready),
    .io_deq_valid(Queue_31_io_deq_valid),
    .io_deq_bits(Queue_31_io_deq_bits)
  );
  assign _T_224_0 = Queue_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18815.4]
  assign _T_224_1 = Queue_1_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18816.4]
  assign _GEN_1 = 4'h1 == auto_in_ar_bits_id ? _T_224_1 : _T_224_0; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_2 = Queue_2_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18817.4]
  assign _GEN_2 = 4'h2 == auto_in_ar_bits_id ? _T_224_2 : _GEN_1; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_3 = Queue_3_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18818.4]
  assign _GEN_3 = 4'h3 == auto_in_ar_bits_id ? _T_224_3 : _GEN_2; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_4 = Queue_4_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18819.4]
  assign _GEN_4 = 4'h4 == auto_in_ar_bits_id ? _T_224_4 : _GEN_3; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_5 = Queue_5_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18820.4]
  assign _GEN_5 = 4'h5 == auto_in_ar_bits_id ? _T_224_5 : _GEN_4; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_6 = Queue_6_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18821.4]
  assign _GEN_6 = 4'h6 == auto_in_ar_bits_id ? _T_224_6 : _GEN_5; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_7 = Queue_7_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18822.4]
  assign _GEN_7 = 4'h7 == auto_in_ar_bits_id ? _T_224_7 : _GEN_6; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_8 = Queue_8_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18823.4]
  assign _GEN_8 = 4'h8 == auto_in_ar_bits_id ? _T_224_8 : _GEN_7; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_9 = Queue_9_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18824.4]
  assign _GEN_9 = 4'h9 == auto_in_ar_bits_id ? _T_224_9 : _GEN_8; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_10 = Queue_10_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18825.4]
  assign _GEN_10 = 4'ha == auto_in_ar_bits_id ? _T_224_10 : _GEN_9; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_11 = Queue_11_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18826.4]
  assign _GEN_11 = 4'hb == auto_in_ar_bits_id ? _T_224_11 : _GEN_10; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_12 = Queue_12_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18827.4]
  assign _GEN_12 = 4'hc == auto_in_ar_bits_id ? _T_224_12 : _GEN_11; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_13 = Queue_13_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18828.4]
  assign _GEN_13 = 4'hd == auto_in_ar_bits_id ? _T_224_13 : _GEN_12; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_14 = Queue_14_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18829.4]
  assign _GEN_14 = 4'he == auto_in_ar_bits_id ? _T_224_14 : _GEN_13; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_224_15 = Queue_15_io_enq_ready; // @[UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18813.4 UserYanker.scala 46:25:boom.system.TestHarness.MegaBoomConfig.fir@18830.4]
  assign _GEN_15 = 4'hf == auto_in_ar_bits_id ? _T_224_15 : _GEN_14; // @[UserYanker.scala 47:36:boom.system.TestHarness.MegaBoomConfig.fir@18831.4]
  assign _T_292 = auto_out_r_valid == 1'h0; // @[UserYanker.scala 54:15:boom.system.TestHarness.MegaBoomConfig.fir@18872.4]
  assign _T_249_0 = Queue_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18838.4]
  assign _T_249_1 = Queue_1_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18839.4]
  assign _GEN_17 = 4'h1 == auto_out_r_bits_id ? _T_249_1 : _T_249_0; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_2 = Queue_2_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18840.4]
  assign _GEN_18 = 4'h2 == auto_out_r_bits_id ? _T_249_2 : _GEN_17; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_3 = Queue_3_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18841.4]
  assign _GEN_19 = 4'h3 == auto_out_r_bits_id ? _T_249_3 : _GEN_18; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_4 = Queue_4_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18842.4]
  assign _GEN_20 = 4'h4 == auto_out_r_bits_id ? _T_249_4 : _GEN_19; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_5 = Queue_5_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18843.4]
  assign _GEN_21 = 4'h5 == auto_out_r_bits_id ? _T_249_5 : _GEN_20; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_6 = Queue_6_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18844.4]
  assign _GEN_22 = 4'h6 == auto_out_r_bits_id ? _T_249_6 : _GEN_21; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_7 = Queue_7_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18845.4]
  assign _GEN_23 = 4'h7 == auto_out_r_bits_id ? _T_249_7 : _GEN_22; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_8 = Queue_8_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18846.4]
  assign _GEN_24 = 4'h8 == auto_out_r_bits_id ? _T_249_8 : _GEN_23; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_9 = Queue_9_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18847.4]
  assign _GEN_25 = 4'h9 == auto_out_r_bits_id ? _T_249_9 : _GEN_24; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_10 = Queue_10_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18848.4]
  assign _GEN_26 = 4'ha == auto_out_r_bits_id ? _T_249_10 : _GEN_25; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_11 = Queue_11_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18849.4]
  assign _GEN_27 = 4'hb == auto_out_r_bits_id ? _T_249_11 : _GEN_26; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_12 = Queue_12_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18850.4]
  assign _GEN_28 = 4'hc == auto_out_r_bits_id ? _T_249_12 : _GEN_27; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_13 = Queue_13_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18851.4]
  assign _GEN_29 = 4'hd == auto_out_r_bits_id ? _T_249_13 : _GEN_28; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_14 = Queue_14_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18852.4]
  assign _GEN_30 = 4'he == auto_out_r_bits_id ? _T_249_14 : _GEN_29; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_249_15 = Queue_15_io_deq_valid; // @[UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18836.4 UserYanker.scala 52:24:boom.system.TestHarness.MegaBoomConfig.fir@18853.4]
  assign _GEN_31 = 4'hf == auto_out_r_bits_id ? _T_249_15 : _GEN_30; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_293 = _T_292 | _GEN_31; // @[UserYanker.scala 54:28:boom.system.TestHarness.MegaBoomConfig.fir@18873.4]
  assign _T_295 = _T_293 | reset; // @[UserYanker.scala 54:14:boom.system.TestHarness.MegaBoomConfig.fir@18875.4]
  assign _T_296 = _T_295 == 1'h0; // @[UserYanker.scala 54:14:boom.system.TestHarness.MegaBoomConfig.fir@18876.4]
  assign _T_272_0 = Queue_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18856.4]
  assign _T_272_1 = Queue_1_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18857.4]
  assign _GEN_33 = 4'h1 == auto_out_r_bits_id ? _T_272_1 : _T_272_0; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_2 = Queue_2_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18858.4]
  assign _GEN_34 = 4'h2 == auto_out_r_bits_id ? _T_272_2 : _GEN_33; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_3 = Queue_3_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18859.4]
  assign _GEN_35 = 4'h3 == auto_out_r_bits_id ? _T_272_3 : _GEN_34; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_4 = Queue_4_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18860.4]
  assign _GEN_36 = 4'h4 == auto_out_r_bits_id ? _T_272_4 : _GEN_35; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_5 = Queue_5_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18861.4]
  assign _GEN_37 = 4'h5 == auto_out_r_bits_id ? _T_272_5 : _GEN_36; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_6 = Queue_6_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18862.4]
  assign _GEN_38 = 4'h6 == auto_out_r_bits_id ? _T_272_6 : _GEN_37; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_7 = Queue_7_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18863.4]
  assign _GEN_39 = 4'h7 == auto_out_r_bits_id ? _T_272_7 : _GEN_38; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_8 = Queue_8_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18864.4]
  assign _GEN_40 = 4'h8 == auto_out_r_bits_id ? _T_272_8 : _GEN_39; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_9 = Queue_9_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18865.4]
  assign _GEN_41 = 4'h9 == auto_out_r_bits_id ? _T_272_9 : _GEN_40; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_10 = Queue_10_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18866.4]
  assign _GEN_42 = 4'ha == auto_out_r_bits_id ? _T_272_10 : _GEN_41; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_11 = Queue_11_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18867.4]
  assign _GEN_43 = 4'hb == auto_out_r_bits_id ? _T_272_11 : _GEN_42; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_12 = Queue_12_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18868.4]
  assign _GEN_44 = 4'hc == auto_out_r_bits_id ? _T_272_12 : _GEN_43; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_13 = Queue_13_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18869.4]
  assign _GEN_45 = 4'hd == auto_out_r_bits_id ? _T_272_13 : _GEN_44; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_14 = Queue_14_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18870.4]
  assign _GEN_46 = 4'he == auto_out_r_bits_id ? _T_272_14 : _GEN_45; // @[UserYanker.scala 56:26:boom.system.TestHarness.MegaBoomConfig.fir@18882.4]
  assign _T_272_15 = Queue_15_io_deq_bits; // @[UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18854.4 UserYanker.scala 53:23:boom.system.TestHarness.MegaBoomConfig.fir@18871.4]
  assign _T_298 = 16'h1 << auto_in_ar_bits_id; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@18884.4]
  assign _T_300 = _T_298[0]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18886.4]
  assign _T_301 = _T_298[1]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18887.4]
  assign _T_302 = _T_298[2]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18888.4]
  assign _T_303 = _T_298[3]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18889.4]
  assign _T_304 = _T_298[4]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18890.4]
  assign _T_305 = _T_298[5]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18891.4]
  assign _T_306 = _T_298[6]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18892.4]
  assign _T_307 = _T_298[7]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18893.4]
  assign _T_308 = _T_298[8]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18894.4]
  assign _T_309 = _T_298[9]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18895.4]
  assign _T_310 = _T_298[10]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18896.4]
  assign _T_311 = _T_298[11]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18897.4]
  assign _T_312 = _T_298[12]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18898.4]
  assign _T_313 = _T_298[13]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18899.4]
  assign _T_314 = _T_298[14]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18900.4]
  assign _T_315 = _T_298[15]; // @[UserYanker.scala 58:55:boom.system.TestHarness.MegaBoomConfig.fir@18901.4]
  assign _T_317 = 16'h1 << auto_out_r_bits_id; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@18903.4]
  assign _T_319 = _T_317[0]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18905.4]
  assign _T_320 = _T_317[1]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18906.4]
  assign _T_321 = _T_317[2]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18907.4]
  assign _T_322 = _T_317[3]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18908.4]
  assign _T_323 = _T_317[4]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18909.4]
  assign _T_324 = _T_317[5]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18910.4]
  assign _T_325 = _T_317[6]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18911.4]
  assign _T_326 = _T_317[7]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18912.4]
  assign _T_327 = _T_317[8]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18913.4]
  assign _T_328 = _T_317[9]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18914.4]
  assign _T_329 = _T_317[10]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18915.4]
  assign _T_330 = _T_317[11]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18916.4]
  assign _T_331 = _T_317[12]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18917.4]
  assign _T_332 = _T_317[13]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18918.4]
  assign _T_333 = _T_317[14]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18919.4]
  assign _T_334 = _T_317[15]; // @[UserYanker.scala 59:55:boom.system.TestHarness.MegaBoomConfig.fir@18920.4]
  assign _T_335 = auto_out_r_valid & auto_in_r_ready; // @[UserYanker.scala 61:37:boom.system.TestHarness.MegaBoomConfig.fir@18921.4]
  assign _T_336 = _T_335 & _T_319; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18922.4]
  assign _T_338 = auto_in_ar_valid & auto_out_ar_ready; // @[UserYanker.scala 62:37:boom.system.TestHarness.MegaBoomConfig.fir@18925.4]
  assign _T_341 = _T_335 & _T_320; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18930.4]
  assign _T_346 = _T_335 & _T_321; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18938.4]
  assign _T_351 = _T_335 & _T_322; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18946.4]
  assign _T_356 = _T_335 & _T_323; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18954.4]
  assign _T_361 = _T_335 & _T_324; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18962.4]
  assign _T_366 = _T_335 & _T_325; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18970.4]
  assign _T_371 = _T_335 & _T_326; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18978.4]
  assign _T_376 = _T_335 & _T_327; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18986.4]
  assign _T_381 = _T_335 & _T_328; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@18994.4]
  assign _T_386 = _T_335 & _T_329; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19002.4]
  assign _T_391 = _T_335 & _T_330; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19010.4]
  assign _T_396 = _T_335 & _T_331; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19018.4]
  assign _T_401 = _T_335 & _T_332; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19026.4]
  assign _T_406 = _T_335 & _T_333; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19034.4]
  assign _T_411 = _T_335 & _T_334; // @[UserYanker.scala 61:53:boom.system.TestHarness.MegaBoomConfig.fir@19042.4]
  assign _T_418_0 = Queue_16_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19051.4]
  assign _T_418_1 = Queue_17_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19052.4]
  assign _GEN_49 = 4'h1 == auto_in_aw_bits_id ? _T_418_1 : _T_418_0; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_2 = Queue_18_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19053.4]
  assign _GEN_50 = 4'h2 == auto_in_aw_bits_id ? _T_418_2 : _GEN_49; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_3 = Queue_19_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19054.4]
  assign _GEN_51 = 4'h3 == auto_in_aw_bits_id ? _T_418_3 : _GEN_50; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_4 = Queue_20_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19055.4]
  assign _GEN_52 = 4'h4 == auto_in_aw_bits_id ? _T_418_4 : _GEN_51; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_5 = Queue_21_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19056.4]
  assign _GEN_53 = 4'h5 == auto_in_aw_bits_id ? _T_418_5 : _GEN_52; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_6 = Queue_22_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19057.4]
  assign _GEN_54 = 4'h6 == auto_in_aw_bits_id ? _T_418_6 : _GEN_53; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_7 = Queue_23_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19058.4]
  assign _GEN_55 = 4'h7 == auto_in_aw_bits_id ? _T_418_7 : _GEN_54; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_8 = Queue_24_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19059.4]
  assign _GEN_56 = 4'h8 == auto_in_aw_bits_id ? _T_418_8 : _GEN_55; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_9 = Queue_25_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19060.4]
  assign _GEN_57 = 4'h9 == auto_in_aw_bits_id ? _T_418_9 : _GEN_56; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_10 = Queue_26_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19061.4]
  assign _GEN_58 = 4'ha == auto_in_aw_bits_id ? _T_418_10 : _GEN_57; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_11 = Queue_27_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19062.4]
  assign _GEN_59 = 4'hb == auto_in_aw_bits_id ? _T_418_11 : _GEN_58; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_12 = Queue_28_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19063.4]
  assign _GEN_60 = 4'hc == auto_in_aw_bits_id ? _T_418_12 : _GEN_59; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_13 = Queue_29_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19064.4]
  assign _GEN_61 = 4'hd == auto_in_aw_bits_id ? _T_418_13 : _GEN_60; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_14 = Queue_30_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19065.4]
  assign _GEN_62 = 4'he == auto_in_aw_bits_id ? _T_418_14 : _GEN_61; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_418_15 = Queue_31_io_enq_ready; // @[UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19049.4 UserYanker.scala 67:25:boom.system.TestHarness.MegaBoomConfig.fir@19066.4]
  assign _GEN_63 = 4'hf == auto_in_aw_bits_id ? _T_418_15 : _GEN_62; // @[UserYanker.scala 68:36:boom.system.TestHarness.MegaBoomConfig.fir@19067.4]
  assign _T_486 = auto_out_b_valid == 1'h0; // @[UserYanker.scala 75:15:boom.system.TestHarness.MegaBoomConfig.fir@19108.4]
  assign _T_443_0 = Queue_16_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19074.4]
  assign _T_443_1 = Queue_17_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19075.4]
  assign _GEN_65 = 4'h1 == auto_out_b_bits_id ? _T_443_1 : _T_443_0; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_2 = Queue_18_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19076.4]
  assign _GEN_66 = 4'h2 == auto_out_b_bits_id ? _T_443_2 : _GEN_65; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_3 = Queue_19_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19077.4]
  assign _GEN_67 = 4'h3 == auto_out_b_bits_id ? _T_443_3 : _GEN_66; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_4 = Queue_20_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19078.4]
  assign _GEN_68 = 4'h4 == auto_out_b_bits_id ? _T_443_4 : _GEN_67; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_5 = Queue_21_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19079.4]
  assign _GEN_69 = 4'h5 == auto_out_b_bits_id ? _T_443_5 : _GEN_68; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_6 = Queue_22_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19080.4]
  assign _GEN_70 = 4'h6 == auto_out_b_bits_id ? _T_443_6 : _GEN_69; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_7 = Queue_23_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19081.4]
  assign _GEN_71 = 4'h7 == auto_out_b_bits_id ? _T_443_7 : _GEN_70; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_8 = Queue_24_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19082.4]
  assign _GEN_72 = 4'h8 == auto_out_b_bits_id ? _T_443_8 : _GEN_71; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_9 = Queue_25_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19083.4]
  assign _GEN_73 = 4'h9 == auto_out_b_bits_id ? _T_443_9 : _GEN_72; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_10 = Queue_26_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19084.4]
  assign _GEN_74 = 4'ha == auto_out_b_bits_id ? _T_443_10 : _GEN_73; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_11 = Queue_27_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19085.4]
  assign _GEN_75 = 4'hb == auto_out_b_bits_id ? _T_443_11 : _GEN_74; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_12 = Queue_28_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19086.4]
  assign _GEN_76 = 4'hc == auto_out_b_bits_id ? _T_443_12 : _GEN_75; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_13 = Queue_29_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19087.4]
  assign _GEN_77 = 4'hd == auto_out_b_bits_id ? _T_443_13 : _GEN_76; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_14 = Queue_30_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19088.4]
  assign _GEN_78 = 4'he == auto_out_b_bits_id ? _T_443_14 : _GEN_77; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_443_15 = Queue_31_io_deq_valid; // @[UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19072.4 UserYanker.scala 73:24:boom.system.TestHarness.MegaBoomConfig.fir@19089.4]
  assign _GEN_79 = 4'hf == auto_out_b_bits_id ? _T_443_15 : _GEN_78; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_487 = _T_486 | _GEN_79; // @[UserYanker.scala 75:28:boom.system.TestHarness.MegaBoomConfig.fir@19109.4]
  assign _T_489 = _T_487 | reset; // @[UserYanker.scala 75:14:boom.system.TestHarness.MegaBoomConfig.fir@19111.4]
  assign _T_490 = _T_489 == 1'h0; // @[UserYanker.scala 75:14:boom.system.TestHarness.MegaBoomConfig.fir@19112.4]
  assign _T_466_0 = Queue_16_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19092.4]
  assign _T_466_1 = Queue_17_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19093.4]
  assign _GEN_81 = 4'h1 == auto_out_b_bits_id ? _T_466_1 : _T_466_0; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_2 = Queue_18_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19094.4]
  assign _GEN_82 = 4'h2 == auto_out_b_bits_id ? _T_466_2 : _GEN_81; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_3 = Queue_19_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19095.4]
  assign _GEN_83 = 4'h3 == auto_out_b_bits_id ? _T_466_3 : _GEN_82; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_4 = Queue_20_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19096.4]
  assign _GEN_84 = 4'h4 == auto_out_b_bits_id ? _T_466_4 : _GEN_83; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_5 = Queue_21_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19097.4]
  assign _GEN_85 = 4'h5 == auto_out_b_bits_id ? _T_466_5 : _GEN_84; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_6 = Queue_22_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19098.4]
  assign _GEN_86 = 4'h6 == auto_out_b_bits_id ? _T_466_6 : _GEN_85; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_7 = Queue_23_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19099.4]
  assign _GEN_87 = 4'h7 == auto_out_b_bits_id ? _T_466_7 : _GEN_86; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_8 = Queue_24_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19100.4]
  assign _GEN_88 = 4'h8 == auto_out_b_bits_id ? _T_466_8 : _GEN_87; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_9 = Queue_25_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19101.4]
  assign _GEN_89 = 4'h9 == auto_out_b_bits_id ? _T_466_9 : _GEN_88; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_10 = Queue_26_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19102.4]
  assign _GEN_90 = 4'ha == auto_out_b_bits_id ? _T_466_10 : _GEN_89; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_11 = Queue_27_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19103.4]
  assign _GEN_91 = 4'hb == auto_out_b_bits_id ? _T_466_11 : _GEN_90; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_12 = Queue_28_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19104.4]
  assign _GEN_92 = 4'hc == auto_out_b_bits_id ? _T_466_12 : _GEN_91; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_13 = Queue_29_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19105.4]
  assign _GEN_93 = 4'hd == auto_out_b_bits_id ? _T_466_13 : _GEN_92; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_14 = Queue_30_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19106.4]
  assign _GEN_94 = 4'he == auto_out_b_bits_id ? _T_466_14 : _GEN_93; // @[UserYanker.scala 77:26:boom.system.TestHarness.MegaBoomConfig.fir@19118.4]
  assign _T_466_15 = Queue_31_io_deq_bits; // @[UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19090.4 UserYanker.scala 74:23:boom.system.TestHarness.MegaBoomConfig.fir@19107.4]
  assign _T_492 = 16'h1 << auto_in_aw_bits_id; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@19120.4]
  assign _T_494 = _T_492[0]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19122.4]
  assign _T_495 = _T_492[1]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19123.4]
  assign _T_496 = _T_492[2]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19124.4]
  assign _T_497 = _T_492[3]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19125.4]
  assign _T_498 = _T_492[4]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19126.4]
  assign _T_499 = _T_492[5]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19127.4]
  assign _T_500 = _T_492[6]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19128.4]
  assign _T_501 = _T_492[7]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19129.4]
  assign _T_502 = _T_492[8]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19130.4]
  assign _T_503 = _T_492[9]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19131.4]
  assign _T_504 = _T_492[10]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19132.4]
  assign _T_505 = _T_492[11]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19133.4]
  assign _T_506 = _T_492[12]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19134.4]
  assign _T_507 = _T_492[13]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19135.4]
  assign _T_508 = _T_492[14]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19136.4]
  assign _T_509 = _T_492[15]; // @[UserYanker.scala 79:55:boom.system.TestHarness.MegaBoomConfig.fir@19137.4]
  assign _T_511 = 16'h1 << auto_out_b_bits_id; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@19139.4]
  assign _T_513 = _T_511[0]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19141.4]
  assign _T_514 = _T_511[1]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19142.4]
  assign _T_515 = _T_511[2]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19143.4]
  assign _T_516 = _T_511[3]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19144.4]
  assign _T_517 = _T_511[4]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19145.4]
  assign _T_518 = _T_511[5]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19146.4]
  assign _T_519 = _T_511[6]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19147.4]
  assign _T_520 = _T_511[7]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19148.4]
  assign _T_521 = _T_511[8]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19149.4]
  assign _T_522 = _T_511[9]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19150.4]
  assign _T_523 = _T_511[10]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19151.4]
  assign _T_524 = _T_511[11]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19152.4]
  assign _T_525 = _T_511[12]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19153.4]
  assign _T_526 = _T_511[13]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19154.4]
  assign _T_527 = _T_511[14]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19155.4]
  assign _T_528 = _T_511[15]; // @[UserYanker.scala 80:55:boom.system.TestHarness.MegaBoomConfig.fir@19156.4]
  assign _T_529 = auto_out_b_valid & auto_in_b_ready; // @[UserYanker.scala 82:37:boom.system.TestHarness.MegaBoomConfig.fir@19157.4]
  assign _T_531 = auto_in_aw_valid & auto_out_aw_ready; // @[UserYanker.scala 83:37:boom.system.TestHarness.MegaBoomConfig.fir@19160.4]
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_63; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_b_bits_user = 4'hf == auto_out_b_bits_id ? _T_466_15 : _GEN_94; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_15; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_r_bits_user = 4'hf == auto_out_r_bits_id ? _T_272_15 : _GEN_46; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@18684.4]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_63; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_15; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@18683.4]
  assign Queue_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18687.4]
  assign Queue_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18688.4]
  assign Queue_io_enq_valid = _T_338 & _T_300; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18927.4]
  assign Queue_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18928.4]
  assign Queue_io_deq_ready = _T_336 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18924.4]
  assign Queue_1_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18691.4]
  assign Queue_1_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18692.4]
  assign Queue_1_io_enq_valid = _T_338 & _T_301; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18935.4]
  assign Queue_1_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18936.4]
  assign Queue_1_io_deq_ready = _T_341 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18932.4]
  assign Queue_2_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18695.4]
  assign Queue_2_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18696.4]
  assign Queue_2_io_enq_valid = _T_338 & _T_302; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18943.4]
  assign Queue_2_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18944.4]
  assign Queue_2_io_deq_ready = _T_346 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18940.4]
  assign Queue_3_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18699.4]
  assign Queue_3_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18700.4]
  assign Queue_3_io_enq_valid = _T_338 & _T_303; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18951.4]
  assign Queue_3_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18952.4]
  assign Queue_3_io_deq_ready = _T_351 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18948.4]
  assign Queue_4_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18703.4]
  assign Queue_4_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18704.4]
  assign Queue_4_io_enq_valid = _T_338 & _T_304; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18959.4]
  assign Queue_4_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18960.4]
  assign Queue_4_io_deq_ready = _T_356 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18956.4]
  assign Queue_5_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18707.4]
  assign Queue_5_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18708.4]
  assign Queue_5_io_enq_valid = _T_338 & _T_305; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18967.4]
  assign Queue_5_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18968.4]
  assign Queue_5_io_deq_ready = _T_361 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18964.4]
  assign Queue_6_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18711.4]
  assign Queue_6_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18712.4]
  assign Queue_6_io_enq_valid = _T_338 & _T_306; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18975.4]
  assign Queue_6_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18976.4]
  assign Queue_6_io_deq_ready = _T_366 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18972.4]
  assign Queue_7_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18715.4]
  assign Queue_7_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18716.4]
  assign Queue_7_io_enq_valid = _T_338 & _T_307; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18983.4]
  assign Queue_7_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18984.4]
  assign Queue_7_io_deq_ready = _T_371 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18980.4]
  assign Queue_8_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18719.4]
  assign Queue_8_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18720.4]
  assign Queue_8_io_enq_valid = _T_338 & _T_308; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18991.4]
  assign Queue_8_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@18992.4]
  assign Queue_8_io_deq_ready = _T_376 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18988.4]
  assign Queue_9_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18723.4]
  assign Queue_9_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18724.4]
  assign Queue_9_io_enq_valid = _T_338 & _T_309; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@18999.4]
  assign Queue_9_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@19000.4]
  assign Queue_9_io_deq_ready = _T_381 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@18996.4]
  assign Queue_10_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18727.4]
  assign Queue_10_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18728.4]
  assign Queue_10_io_enq_valid = _T_338 & _T_310; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@19007.4]
  assign Queue_10_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@19008.4]
  assign Queue_10_io_deq_ready = _T_386 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@19004.4]
  assign Queue_11_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18731.4]
  assign Queue_11_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18732.4]
  assign Queue_11_io_enq_valid = _T_338 & _T_311; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@19015.4]
  assign Queue_11_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@19016.4]
  assign Queue_11_io_deq_ready = _T_391 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@19012.4]
  assign Queue_12_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18735.4]
  assign Queue_12_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18736.4]
  assign Queue_12_io_enq_valid = _T_338 & _T_312; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@19023.4]
  assign Queue_12_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@19024.4]
  assign Queue_12_io_deq_ready = _T_396 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@19020.4]
  assign Queue_13_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18739.4]
  assign Queue_13_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18740.4]
  assign Queue_13_io_enq_valid = _T_338 & _T_313; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@19031.4]
  assign Queue_13_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@19032.4]
  assign Queue_13_io_deq_ready = _T_401 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@19028.4]
  assign Queue_14_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18743.4]
  assign Queue_14_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18744.4]
  assign Queue_14_io_enq_valid = _T_338 & _T_314; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@19039.4]
  assign Queue_14_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@19040.4]
  assign Queue_14_io_deq_ready = _T_406 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@19036.4]
  assign Queue_15_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18747.4]
  assign Queue_15_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18748.4]
  assign Queue_15_io_enq_valid = _T_338 & _T_315; // @[UserYanker.scala 62:21:boom.system.TestHarness.MegaBoomConfig.fir@19047.4]
  assign Queue_15_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:boom.system.TestHarness.MegaBoomConfig.fir@19048.4]
  assign Queue_15_io_deq_ready = _T_411 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:boom.system.TestHarness.MegaBoomConfig.fir@19044.4]
  assign Queue_16_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18751.4]
  assign Queue_16_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18752.4]
  assign Queue_16_io_enq_valid = _T_531 & _T_494; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19162.4]
  assign Queue_16_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19163.4]
  assign Queue_16_io_deq_ready = _T_529 & _T_513; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19159.4]
  assign Queue_17_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18755.4]
  assign Queue_17_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18756.4]
  assign Queue_17_io_enq_valid = _T_531 & _T_495; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19169.4]
  assign Queue_17_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19170.4]
  assign Queue_17_io_deq_ready = _T_529 & _T_514; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19166.4]
  assign Queue_18_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18759.4]
  assign Queue_18_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18760.4]
  assign Queue_18_io_enq_valid = _T_531 & _T_496; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19176.4]
  assign Queue_18_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19177.4]
  assign Queue_18_io_deq_ready = _T_529 & _T_515; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19173.4]
  assign Queue_19_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18763.4]
  assign Queue_19_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18764.4]
  assign Queue_19_io_enq_valid = _T_531 & _T_497; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19183.4]
  assign Queue_19_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19184.4]
  assign Queue_19_io_deq_ready = _T_529 & _T_516; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19180.4]
  assign Queue_20_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18767.4]
  assign Queue_20_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18768.4]
  assign Queue_20_io_enq_valid = _T_531 & _T_498; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19190.4]
  assign Queue_20_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19191.4]
  assign Queue_20_io_deq_ready = _T_529 & _T_517; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19187.4]
  assign Queue_21_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18771.4]
  assign Queue_21_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18772.4]
  assign Queue_21_io_enq_valid = _T_531 & _T_499; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19197.4]
  assign Queue_21_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19198.4]
  assign Queue_21_io_deq_ready = _T_529 & _T_518; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19194.4]
  assign Queue_22_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18775.4]
  assign Queue_22_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18776.4]
  assign Queue_22_io_enq_valid = _T_531 & _T_500; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19204.4]
  assign Queue_22_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19205.4]
  assign Queue_22_io_deq_ready = _T_529 & _T_519; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19201.4]
  assign Queue_23_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18779.4]
  assign Queue_23_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18780.4]
  assign Queue_23_io_enq_valid = _T_531 & _T_501; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19211.4]
  assign Queue_23_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19212.4]
  assign Queue_23_io_deq_ready = _T_529 & _T_520; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19208.4]
  assign Queue_24_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18783.4]
  assign Queue_24_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18784.4]
  assign Queue_24_io_enq_valid = _T_531 & _T_502; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19218.4]
  assign Queue_24_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19219.4]
  assign Queue_24_io_deq_ready = _T_529 & _T_521; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19215.4]
  assign Queue_25_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18787.4]
  assign Queue_25_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18788.4]
  assign Queue_25_io_enq_valid = _T_531 & _T_503; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19225.4]
  assign Queue_25_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19226.4]
  assign Queue_25_io_deq_ready = _T_529 & _T_522; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19222.4]
  assign Queue_26_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18791.4]
  assign Queue_26_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18792.4]
  assign Queue_26_io_enq_valid = _T_531 & _T_504; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19232.4]
  assign Queue_26_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19233.4]
  assign Queue_26_io_deq_ready = _T_529 & _T_523; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19229.4]
  assign Queue_27_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18795.4]
  assign Queue_27_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18796.4]
  assign Queue_27_io_enq_valid = _T_531 & _T_505; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19239.4]
  assign Queue_27_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19240.4]
  assign Queue_27_io_deq_ready = _T_529 & _T_524; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19236.4]
  assign Queue_28_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18799.4]
  assign Queue_28_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18800.4]
  assign Queue_28_io_enq_valid = _T_531 & _T_506; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19246.4]
  assign Queue_28_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19247.4]
  assign Queue_28_io_deq_ready = _T_529 & _T_525; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19243.4]
  assign Queue_29_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18803.4]
  assign Queue_29_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18804.4]
  assign Queue_29_io_enq_valid = _T_531 & _T_507; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19253.4]
  assign Queue_29_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19254.4]
  assign Queue_29_io_deq_ready = _T_529 & _T_526; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19250.4]
  assign Queue_30_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18807.4]
  assign Queue_30_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18808.4]
  assign Queue_30_io_enq_valid = _T_531 & _T_508; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19260.4]
  assign Queue_30_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19261.4]
  assign Queue_30_io_deq_ready = _T_529 & _T_527; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19257.4]
  assign Queue_31_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18811.4]
  assign Queue_31_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@18812.4]
  assign Queue_31_io_enq_valid = _T_531 & _T_509; // @[UserYanker.scala 83:21:boom.system.TestHarness.MegaBoomConfig.fir@19267.4]
  assign Queue_31_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:boom.system.TestHarness.MegaBoomConfig.fir@19268.4]
  assign Queue_31_io_deq_ready = _T_529 & _T_528; // @[UserYanker.scala 82:21:boom.system.TestHarness.MegaBoomConfig.fir@19264.4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_296) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:54 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"); // @[UserYanker.scala 54:14:boom.system.TestHarness.MegaBoomConfig.fir@18878.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_296) begin
          $fatal; // @[UserYanker.scala 54:14:boom.system.TestHarness.MegaBoomConfig.fir@18879.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_490) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:75 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"); // @[UserYanker.scala 75:14:boom.system.TestHarness.MegaBoomConfig.fir@19114.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_490) begin
          $fatal; // @[UserYanker.scala 75:14:boom.system.TestHarness.MegaBoomConfig.fir@19115.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer_2( // @[:boom.system.TestHarness.MegaBoomConfig.fir@19271.2]
  output        auto_in_aw_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_in_aw_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [7:0]  auto_in_aw_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [31:0] auto_in_aw_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_in_aw_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [11:0] auto_in_aw_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_in_w_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_in_w_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [63:0] auto_in_w_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [7:0]  auto_in_w_bits_strb, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_in_w_bits_last, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_in_b_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_in_b_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [7:0]  auto_in_b_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [1:0]  auto_in_b_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [11:0] auto_in_b_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_in_ar_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_in_ar_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [7:0]  auto_in_ar_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [31:0] auto_in_ar_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_in_ar_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [11:0] auto_in_ar_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_in_r_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_in_r_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [7:0]  auto_in_r_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [63:0] auto_in_r_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [1:0]  auto_in_r_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [11:0] auto_in_r_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_in_r_bits_last, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_out_aw_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_out_aw_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [3:0]  auto_out_aw_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [31:0] auto_out_aw_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [7:0]  auto_out_aw_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [2:0]  auto_out_aw_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_out_aw_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [15:0] auto_out_aw_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_out_w_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_out_w_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [63:0] auto_out_w_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [7:0]  auto_out_w_bits_strb, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_out_w_bits_last, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_out_b_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_out_b_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [3:0]  auto_out_b_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [15:0] auto_out_b_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_out_ar_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_out_ar_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [3:0]  auto_out_ar_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [31:0] auto_out_ar_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [7:0]  auto_out_ar_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [2:0]  auto_out_ar_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_out_ar_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output [15:0] auto_out_ar_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  output        auto_out_r_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_out_r_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [3:0]  auto_out_r_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [63:0] auto_out_r_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input  [15:0] auto_out_r_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
  input         auto_out_r_bits_last // @[:boom.system.TestHarness.MegaBoomConfig.fir@19274.4]
);
  wire [3:0] _T_221; // @[IdIndexer.scala 56:81:boom.system.TestHarness.MegaBoomConfig.fir@19290.4]
  wire [3:0] _T_223; // @[IdIndexer.scala 57:81:boom.system.TestHarness.MegaBoomConfig.fir@19293.4]
  wire [19:0] _T_227; // @[Cat.scala 30:58:boom.system.TestHarness.MegaBoomConfig.fir@19300.4]
  wire [19:0] _T_228; // @[Cat.scala 30:58:boom.system.TestHarness.MegaBoomConfig.fir@19302.4]
  assign _T_221 = auto_in_ar_bits_id[7:4]; // @[IdIndexer.scala 56:81:boom.system.TestHarness.MegaBoomConfig.fir@19290.4]
  assign _T_223 = auto_in_aw_bits_id[7:4]; // @[IdIndexer.scala 57:81:boom.system.TestHarness.MegaBoomConfig.fir@19293.4]
  assign _T_227 = {auto_out_r_bits_user,auto_out_r_bits_id}; // @[Cat.scala 30:58:boom.system.TestHarness.MegaBoomConfig.fir@19300.4]
  assign _T_228 = {auto_out_b_bits_user,auto_out_b_bits_id}; // @[Cat.scala 30:58:boom.system.TestHarness.MegaBoomConfig.fir@19302.4]
  assign auto_in_aw_ready = auto_out_aw_ready; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_b_bits_id = _T_228[7:0]; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_b_bits_user = auto_out_b_bits_user[15:4]; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_r_bits_id = _T_227[7:0]; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_r_bits_user = auto_out_r_bits_user[15:4]; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19284.4]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id[3:0]; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_aw_bits_user = {auto_in_aw_bits_user,_T_223}; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id[3:0]; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_ar_bits_user = {auto_in_ar_bits_user,_T_221}; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19283.4]
endmodule
module Queue_97( // @[:boom.system.TestHarness.MegaBoomConfig.fir@19361.2]
  input         clock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19362.4]
  input         reset, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19363.4]
  output        io_enq_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  input         io_enq_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  input  [7:0]  io_enq_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  input  [31:0] io_enq_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  input  [7:0]  io_enq_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  input  [2:0]  io_enq_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  input  [11:0] io_enq_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  input         io_enq_bits_wen, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  input         io_deq_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output        io_deq_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [7:0]  io_deq_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [31:0] io_deq_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [7:0]  io_deq_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [2:0]  io_deq_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [1:0]  io_deq_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output        io_deq_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [3:0]  io_deq_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [2:0]  io_deq_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [3:0]  io_deq_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output [11:0] io_deq_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
  output        io_deq_bits_wen // @[:boom.system.TestHarness.MegaBoomConfig.fir@19364.4]
);
  reg [7:0] _T_35_id [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_0;
  wire [7:0] _T_35_id__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_id__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [7:0] _T_35_id__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_id__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_id__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_id__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _T_35_addr [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_1;
  wire [31:0] _T_35_addr__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_addr__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [31:0] _T_35_addr__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_addr__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_addr__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_addr__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [7:0] _T_35_len [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_2;
  wire [7:0] _T_35_len__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_len__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [7:0] _T_35_len__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_len__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_len__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_len__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [2:0] _T_35_size [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_3;
  wire [2:0] _T_35_size__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_size__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [2:0] _T_35_size__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_size__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_size__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_size__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [1:0] _T_35_burst [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_4;
  wire [1:0] _T_35_burst__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_burst__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [1:0] _T_35_burst__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_burst__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_burst__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_burst__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg  _T_35_lock [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_5;
  wire  _T_35_lock__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_lock__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_lock__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_lock__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_lock__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_lock__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [3:0] _T_35_cache [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_6;
  wire [3:0] _T_35_cache__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_cache__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [3:0] _T_35_cache__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_cache__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_cache__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_cache__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [2:0] _T_35_prot [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_7;
  wire [2:0] _T_35_prot__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_prot__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [2:0] _T_35_prot__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_prot__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_prot__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_prot__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [3:0] _T_35_qos [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_8;
  wire [3:0] _T_35_qos__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_qos__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [3:0] _T_35_qos__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_qos__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_qos__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_qos__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [11:0] _T_35_user [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_9;
  wire [11:0] _T_35_user__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_user__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire [11:0] _T_35_user__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_user__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_user__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_user__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg  _T_35_wen [0:0]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg [31:0] _RAND_10;
  wire  _T_35_wen__T_52_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_wen__T_52_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_wen__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_wen__T_48_addr; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_wen__T_48_mask; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  wire  _T_35_wen__T_48_en; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  reg  _T_37; // @[Decoupled.scala 217:35:boom.system.TestHarness.MegaBoomConfig.fir@19367.4]
  reg [31:0] _RAND_11;
  wire  _T_39; // @[Decoupled.scala 220:36:boom.system.TestHarness.MegaBoomConfig.fir@19369.4]
  wire  _T_42; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@19372.4]
  wire  _T_45; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@19375.4]
  wire  _GEN_17; // @[Decoupled.scala 245:27:boom.system.TestHarness.MegaBoomConfig.fir@19430.6]
  wire  _GEN_30; // @[Decoupled.scala 242:18:boom.system.TestHarness.MegaBoomConfig.fir@19417.4]
  wire  _GEN_29; // @[Decoupled.scala 242:18:boom.system.TestHarness.MegaBoomConfig.fir@19417.4]
  wire  _T_49; // @[Decoupled.scala 232:16:boom.system.TestHarness.MegaBoomConfig.fir@19394.4]
  wire  _T_50; // @[Decoupled.scala 236:19:boom.system.TestHarness.MegaBoomConfig.fir@19398.4]
  assign _T_35_id__T_52_addr = 1'h0;
  assign _T_35_id__T_52_data = _T_35_id[_T_35_id__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_id__T_48_data = io_enq_bits_id;
  assign _T_35_id__T_48_addr = 1'h0;
  assign _T_35_id__T_48_mask = 1'h1;
  assign _T_35_id__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_addr__T_52_addr = 1'h0;
  assign _T_35_addr__T_52_data = _T_35_addr[_T_35_addr__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_addr__T_48_data = io_enq_bits_addr;
  assign _T_35_addr__T_48_addr = 1'h0;
  assign _T_35_addr__T_48_mask = 1'h1;
  assign _T_35_addr__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_len__T_52_addr = 1'h0;
  assign _T_35_len__T_52_data = _T_35_len[_T_35_len__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_len__T_48_data = io_enq_bits_len;
  assign _T_35_len__T_48_addr = 1'h0;
  assign _T_35_len__T_48_mask = 1'h1;
  assign _T_35_len__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_size__T_52_addr = 1'h0;
  assign _T_35_size__T_52_data = _T_35_size[_T_35_size__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_size__T_48_data = io_enq_bits_size;
  assign _T_35_size__T_48_addr = 1'h0;
  assign _T_35_size__T_48_mask = 1'h1;
  assign _T_35_size__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_burst__T_52_addr = 1'h0;
  assign _T_35_burst__T_52_data = _T_35_burst[_T_35_burst__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_burst__T_48_data = 2'h1;
  assign _T_35_burst__T_48_addr = 1'h0;
  assign _T_35_burst__T_48_mask = 1'h1;
  assign _T_35_burst__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_lock__T_52_addr = 1'h0;
  assign _T_35_lock__T_52_data = _T_35_lock[_T_35_lock__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_lock__T_48_data = 1'h0;
  assign _T_35_lock__T_48_addr = 1'h0;
  assign _T_35_lock__T_48_mask = 1'h1;
  assign _T_35_lock__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_cache__T_52_addr = 1'h0;
  assign _T_35_cache__T_52_data = _T_35_cache[_T_35_cache__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_cache__T_48_data = 4'h0;
  assign _T_35_cache__T_48_addr = 1'h0;
  assign _T_35_cache__T_48_mask = 1'h1;
  assign _T_35_cache__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_prot__T_52_addr = 1'h0;
  assign _T_35_prot__T_52_data = _T_35_prot[_T_35_prot__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_prot__T_48_data = 3'h1;
  assign _T_35_prot__T_48_addr = 1'h0;
  assign _T_35_prot__T_48_mask = 1'h1;
  assign _T_35_prot__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_qos__T_52_addr = 1'h0;
  assign _T_35_qos__T_52_data = _T_35_qos[_T_35_qos__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_qos__T_48_data = 4'h0;
  assign _T_35_qos__T_48_addr = 1'h0;
  assign _T_35_qos__T_48_mask = 1'h1;
  assign _T_35_qos__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_user__T_52_addr = 1'h0;
  assign _T_35_user__T_52_data = _T_35_user[_T_35_user__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_user__T_48_data = io_enq_bits_user;
  assign _T_35_user__T_48_addr = 1'h0;
  assign _T_35_user__T_48_mask = 1'h1;
  assign _T_35_user__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_wen__T_52_addr = 1'h0;
  assign _T_35_wen__T_52_data = _T_35_wen[_T_35_wen__T_52_addr]; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
  assign _T_35_wen__T_48_data = io_enq_bits_wen;
  assign _T_35_wen__T_48_addr = 1'h0;
  assign _T_35_wen__T_48_mask = 1'h1;
  assign _T_35_wen__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_39 = _T_37 == 1'h0; // @[Decoupled.scala 220:36:boom.system.TestHarness.MegaBoomConfig.fir@19369.4]
  assign _T_42 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@19372.4]
  assign _T_45 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@19375.4]
  assign _GEN_17 = io_deq_ready ? 1'h0 : _T_42; // @[Decoupled.scala 245:27:boom.system.TestHarness.MegaBoomConfig.fir@19430.6]
  assign _GEN_30 = _T_39 ? _GEN_17 : _T_42; // @[Decoupled.scala 242:18:boom.system.TestHarness.MegaBoomConfig.fir@19417.4]
  assign _GEN_29 = _T_39 ? 1'h0 : _T_45; // @[Decoupled.scala 242:18:boom.system.TestHarness.MegaBoomConfig.fir@19417.4]
  assign _T_49 = _GEN_30 != _GEN_29; // @[Decoupled.scala 232:16:boom.system.TestHarness.MegaBoomConfig.fir@19394.4]
  assign _T_50 = _T_39 == 1'h0; // @[Decoupled.scala 236:19:boom.system.TestHarness.MegaBoomConfig.fir@19398.4]
  assign io_enq_ready = _T_37 == 1'h0; // @[Decoupled.scala 237:16:boom.system.TestHarness.MegaBoomConfig.fir@19401.4]
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_50; // @[Decoupled.scala 236:16:boom.system.TestHarness.MegaBoomConfig.fir@19399.4 Decoupled.scala 241:40:boom.system.TestHarness.MegaBoomConfig.fir@19415.6]
  assign io_deq_bits_id = _T_39 ? io_enq_bits_id : _T_35_id__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19413.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19428.6]
  assign io_deq_bits_addr = _T_39 ? io_enq_bits_addr : _T_35_addr__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19412.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19427.6]
  assign io_deq_bits_len = _T_39 ? io_enq_bits_len : _T_35_len__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19411.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19426.6]
  assign io_deq_bits_size = _T_39 ? io_enq_bits_size : _T_35_size__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19410.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19425.6]
  assign io_deq_bits_burst = _T_39 ? 2'h1 : _T_35_burst__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19409.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19424.6]
  assign io_deq_bits_lock = _T_39 ? 1'h0 : _T_35_lock__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19408.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19423.6]
  assign io_deq_bits_cache = _T_39 ? 4'h0 : _T_35_cache__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19407.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19422.6]
  assign io_deq_bits_prot = _T_39 ? 3'h1 : _T_35_prot__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19406.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19421.6]
  assign io_deq_bits_qos = _T_39 ? 4'h0 : _T_35_qos__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19405.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19420.6]
  assign io_deq_bits_user = _T_39 ? io_enq_bits_user : _T_35_user__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19404.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19419.6]
  assign io_deq_bits_wen = _T_39 ? io_enq_bits_wen : _T_35_wen__T_52_data; // @[Decoupled.scala 238:15:boom.system.TestHarness.MegaBoomConfig.fir@19403.4 Decoupled.scala 243:19:boom.system.TestHarness.MegaBoomConfig.fir@19418.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_id[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_addr[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_user[initvar] = _RAND_9[11:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_wen[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_37 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35_id__T_48_en & _T_35_id__T_48_mask) begin
      _T_35_id[_T_35_id__T_48_addr] <= _T_35_id__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_addr__T_48_en & _T_35_addr__T_48_mask) begin
      _T_35_addr[_T_35_addr__T_48_addr] <= _T_35_addr__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_len__T_48_en & _T_35_len__T_48_mask) begin
      _T_35_len[_T_35_len__T_48_addr] <= _T_35_len__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_size__T_48_en & _T_35_size__T_48_mask) begin
      _T_35_size[_T_35_size__T_48_addr] <= _T_35_size__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_burst__T_48_en & _T_35_burst__T_48_mask) begin
      _T_35_burst[_T_35_burst__T_48_addr] <= _T_35_burst__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_lock__T_48_en & _T_35_lock__T_48_mask) begin
      _T_35_lock[_T_35_lock__T_48_addr] <= _T_35_lock__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_cache__T_48_en & _T_35_cache__T_48_mask) begin
      _T_35_cache[_T_35_cache__T_48_addr] <= _T_35_cache__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_prot__T_48_en & _T_35_prot__T_48_mask) begin
      _T_35_prot[_T_35_prot__T_48_addr] <= _T_35_prot__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_qos__T_48_en & _T_35_qos__T_48_mask) begin
      _T_35_qos[_T_35_qos__T_48_addr] <= _T_35_qos__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_user__T_48_en & _T_35_user__T_48_mask) begin
      _T_35_user[_T_35_user__T_48_addr] <= _T_35_user__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if(_T_35_wen__T_48_en & _T_35_wen__T_48_mask) begin
      _T_35_wen[_T_35_wen__T_48_addr] <= _T_35_wen__T_48_data; // @[Decoupled.scala 214:24:boom.system.TestHarness.MegaBoomConfig.fir@19366.4]
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_49) begin
        if (_T_39) begin
          if (io_deq_ready) begin
            _T_37 <= 1'h0;
          end else begin
            _T_37 <= _T_42;
          end
        end else begin
          _T_37 <= _T_42;
        end
      end
    end
  end
endmodule
module TLToAXI4_1( // @[:boom.system.TestHarness.MegaBoomConfig.fir@19441.2]
  input         clock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19442.4]
  input         reset, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19443.4]
  output        auto_in_a_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input         auto_in_a_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [2:0]  auto_in_a_bits_opcode, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [2:0]  auto_in_a_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [7:0]  auto_in_a_bits_source, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [31:0] auto_in_a_bits_address, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [7:0]  auto_in_a_bits_mask, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [63:0] auto_in_a_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input         auto_in_d_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_in_d_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [2:0]  auto_in_d_bits_opcode, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [2:0]  auto_in_d_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [7:0]  auto_in_d_bits_source, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_in_d_bits_denied, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [63:0] auto_in_d_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_in_d_bits_corrupt, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input         auto_out_aw_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_out_aw_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [7:0]  auto_out_aw_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [31:0] auto_out_aw_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [7:0]  auto_out_aw_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [2:0]  auto_out_aw_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_out_aw_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [11:0] auto_out_aw_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input         auto_out_w_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_out_w_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [63:0] auto_out_w_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [7:0]  auto_out_w_bits_strb, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_out_w_bits_last, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_out_b_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input         auto_out_b_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [7:0]  auto_out_b_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [11:0] auto_out_b_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input         auto_out_ar_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_out_ar_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [7:0]  auto_out_ar_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [31:0] auto_out_ar_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [7:0]  auto_out_ar_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [2:0]  auto_out_ar_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_out_ar_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output [11:0] auto_out_ar_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  output        auto_out_r_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input         auto_out_r_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [7:0]  auto_out_r_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [63:0] auto_out_r_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input  [11:0] auto_out_r_bits_user, // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
  input         auto_out_r_bits_last // @[:boom.system.TestHarness.MegaBoomConfig.fir@19444.4]
);
  wire  Queue_clock; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire  Queue_reset; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire [63:0] Queue_io_enq_bits_data; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire [7:0] Queue_io_enq_bits_strb; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire [63:0] Queue_io_deq_bits_data; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire [7:0] Queue_io_deq_bits_strb; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
  wire  Queue_1_clock; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  Queue_1_reset; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [7:0] Queue_1_io_enq_bits_id; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [31:0] Queue_1_io_enq_bits_addr; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [7:0] Queue_1_io_enq_bits_len; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [2:0] Queue_1_io_enq_bits_size; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [11:0] Queue_1_io_enq_bits_user; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  Queue_1_io_enq_bits_wen; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [7:0] Queue_1_io_deq_bits_id; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [31:0] Queue_1_io_deq_bits_addr; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [7:0] Queue_1_io_deq_bits_len; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [2:0] Queue_1_io_deq_bits_size; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [1:0] Queue_1_io_deq_bits_burst; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  Queue_1_io_deq_bits_lock; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [3:0] Queue_1_io_deq_bits_cache; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [2:0] Queue_1_io_deq_bits_prot; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [3:0] Queue_1_io_deq_bits_qos; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire [11:0] Queue_1_io_deq_bits_user; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  Queue_1_io_deq_bits_wen; // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
  wire  _T_2295; // @[Edges.scala 92:37:boom.system.TestHarness.MegaBoomConfig.fir@20232.4]
  wire  _T_2296; // @[Edges.scala 92:28:boom.system.TestHarness.MegaBoomConfig.fir@20233.4]
  reg  _T_10843; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31666.4]
  reg [31:0] _RAND_0;
  reg  _T_10812; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31624.4]
  reg [31:0] _RAND_1;
  reg  _T_10781; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31582.4]
  reg [31:0] _RAND_2;
  reg  _T_10750; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31540.4]
  reg [31:0] _RAND_3;
  reg  _T_10719; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31498.4]
  reg [31:0] _RAND_4;
  reg  _T_10688; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31456.4]
  reg [31:0] _RAND_5;
  reg  _T_10657; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31414.4]
  reg [31:0] _RAND_6;
  reg  _T_10626; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31372.4]
  reg [31:0] _RAND_7;
  reg  _T_10595; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31330.4]
  reg [31:0] _RAND_8;
  reg  _T_10564; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31288.4]
  reg [31:0] _RAND_9;
  reg  _T_10533; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31246.4]
  reg [31:0] _RAND_10;
  reg  _T_10502; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31204.4]
  reg [31:0] _RAND_11;
  reg  _T_10471; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31162.4]
  reg [31:0] _RAND_12;
  reg  _T_10440; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31120.4]
  reg [31:0] _RAND_13;
  reg  _T_10409; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31078.4]
  reg [31:0] _RAND_14;
  reg  _T_10378; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@31036.4]
  reg [31:0] _RAND_15;
  reg  _T_10347; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30994.4]
  reg [31:0] _RAND_16;
  reg  _T_10316; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30952.4]
  reg [31:0] _RAND_17;
  reg  _T_10285; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30910.4]
  reg [31:0] _RAND_18;
  reg  _T_10254; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30868.4]
  reg [31:0] _RAND_19;
  reg  _T_10223; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30826.4]
  reg [31:0] _RAND_20;
  reg  _T_10192; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30784.4]
  reg [31:0] _RAND_21;
  reg  _T_10161; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30742.4]
  reg [31:0] _RAND_22;
  reg  _T_10130; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30700.4]
  reg [31:0] _RAND_23;
  reg  _T_10099; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30658.4]
  reg [31:0] _RAND_24;
  reg  _T_10068; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30616.4]
  reg [31:0] _RAND_25;
  reg  _T_10037; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30574.4]
  reg [31:0] _RAND_26;
  reg  _T_10006; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30532.4]
  reg [31:0] _RAND_27;
  reg  _T_9975; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30490.4]
  reg [31:0] _RAND_28;
  reg  _T_9944; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30448.4]
  reg [31:0] _RAND_29;
  reg  _T_9913; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30406.4]
  reg [31:0] _RAND_30;
  reg  _T_9882; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30364.4]
  reg [31:0] _RAND_31;
  reg  _T_9851; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30322.4]
  reg [31:0] _RAND_32;
  reg  _T_9820; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30280.4]
  reg [31:0] _RAND_33;
  reg  _T_9789; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30238.4]
  reg [31:0] _RAND_34;
  reg  _T_9758; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30196.4]
  reg [31:0] _RAND_35;
  reg  _T_9727; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30154.4]
  reg [31:0] _RAND_36;
  reg  _T_9696; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30112.4]
  reg [31:0] _RAND_37;
  reg  _T_9665; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30070.4]
  reg [31:0] _RAND_38;
  reg  _T_9634; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@30028.4]
  reg [31:0] _RAND_39;
  reg  _T_9603; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29986.4]
  reg [31:0] _RAND_40;
  reg  _T_9572; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29944.4]
  reg [31:0] _RAND_41;
  reg  _T_9541; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29902.4]
  reg [31:0] _RAND_42;
  reg  _T_9510; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29860.4]
  reg [31:0] _RAND_43;
  reg  _T_9479; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29818.4]
  reg [31:0] _RAND_44;
  reg  _T_9448; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29776.4]
  reg [31:0] _RAND_45;
  reg  _T_9417; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29734.4]
  reg [31:0] _RAND_46;
  reg  _T_9386; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29692.4]
  reg [31:0] _RAND_47;
  reg  _T_9355; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29650.4]
  reg [31:0] _RAND_48;
  reg  _T_9324; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29608.4]
  reg [31:0] _RAND_49;
  reg  _T_9293; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29566.4]
  reg [31:0] _RAND_50;
  reg  _T_9262; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29524.4]
  reg [31:0] _RAND_51;
  reg  _T_9231; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29482.4]
  reg [31:0] _RAND_52;
  reg  _T_9200; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29440.4]
  reg [31:0] _RAND_53;
  reg  _T_9169; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29398.4]
  reg [31:0] _RAND_54;
  reg  _T_9138; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29356.4]
  reg [31:0] _RAND_55;
  reg  _T_9107; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29314.4]
  reg [31:0] _RAND_56;
  reg  _T_9076; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29272.4]
  reg [31:0] _RAND_57;
  reg  _T_9045; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29230.4]
  reg [31:0] _RAND_58;
  reg  _T_9014; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29188.4]
  reg [31:0] _RAND_59;
  reg  _T_8983; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29146.4]
  reg [31:0] _RAND_60;
  reg  _T_8952; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29104.4]
  reg [31:0] _RAND_61;
  reg  _T_8921; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29062.4]
  reg [31:0] _RAND_62;
  reg  _T_8890; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@29020.4]
  reg [31:0] _RAND_63;
  reg  _T_8859; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28978.4]
  reg [31:0] _RAND_64;
  reg  _T_8828; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28936.4]
  reg [31:0] _RAND_65;
  reg  _T_8797; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28894.4]
  reg [31:0] _RAND_66;
  reg  _T_8766; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28852.4]
  reg [31:0] _RAND_67;
  reg  _T_8735; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28810.4]
  reg [31:0] _RAND_68;
  reg  _T_8704; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28768.4]
  reg [31:0] _RAND_69;
  reg  _T_8673; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28726.4]
  reg [31:0] _RAND_70;
  reg  _T_8642; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28684.4]
  reg [31:0] _RAND_71;
  reg  _T_8611; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28642.4]
  reg [31:0] _RAND_72;
  reg  _T_8580; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28600.4]
  reg [31:0] _RAND_73;
  reg  _T_8549; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28558.4]
  reg [31:0] _RAND_74;
  reg  _T_8518; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28516.4]
  reg [31:0] _RAND_75;
  reg  _T_8487; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28474.4]
  reg [31:0] _RAND_76;
  reg  _T_8456; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28432.4]
  reg [31:0] _RAND_77;
  reg  _T_8425; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28390.4]
  reg [31:0] _RAND_78;
  reg  _T_8394; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28348.4]
  reg [31:0] _RAND_79;
  reg  _T_8363; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28306.4]
  reg [31:0] _RAND_80;
  reg  _T_8332; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28264.4]
  reg [31:0] _RAND_81;
  reg  _T_8301; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28222.4]
  reg [31:0] _RAND_82;
  reg  _T_8270; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28180.4]
  reg [31:0] _RAND_83;
  reg  _T_8239; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28138.4]
  reg [31:0] _RAND_84;
  reg  _T_8208; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28096.4]
  reg [31:0] _RAND_85;
  reg  _T_8177; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28054.4]
  reg [31:0] _RAND_86;
  reg  _T_8146; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@28012.4]
  reg [31:0] _RAND_87;
  reg  _T_8115; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27970.4]
  reg [31:0] _RAND_88;
  reg  _T_8084; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27928.4]
  reg [31:0] _RAND_89;
  reg  _T_8053; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27886.4]
  reg [31:0] _RAND_90;
  reg  _T_8022; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27844.4]
  reg [31:0] _RAND_91;
  reg  _T_7991; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27802.4]
  reg [31:0] _RAND_92;
  reg  _T_7960; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27760.4]
  reg [31:0] _RAND_93;
  reg  _T_7929; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27718.4]
  reg [31:0] _RAND_94;
  reg  _T_7898; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27676.4]
  reg [31:0] _RAND_95;
  reg  _T_7867; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27634.4]
  reg [31:0] _RAND_96;
  reg  _T_7836; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27592.4]
  reg [31:0] _RAND_97;
  reg  _T_7805; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27550.4]
  reg [31:0] _RAND_98;
  reg  _T_7774; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27508.4]
  reg [31:0] _RAND_99;
  reg  _T_7743; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27466.4]
  reg [31:0] _RAND_100;
  reg  _T_7712; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27424.4]
  reg [31:0] _RAND_101;
  reg  _T_7681; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27382.4]
  reg [31:0] _RAND_102;
  reg  _T_7650; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27340.4]
  reg [31:0] _RAND_103;
  reg  _T_7619; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27298.4]
  reg [31:0] _RAND_104;
  reg  _T_7588; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27256.4]
  reg [31:0] _RAND_105;
  reg  _T_7557; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27214.4]
  reg [31:0] _RAND_106;
  reg  _T_7526; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27172.4]
  reg [31:0] _RAND_107;
  reg  _T_7495; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27130.4]
  reg [31:0] _RAND_108;
  reg  _T_7464; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27088.4]
  reg [31:0] _RAND_109;
  reg  _T_7433; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27046.4]
  reg [31:0] _RAND_110;
  reg  _T_7402; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@27004.4]
  reg [31:0] _RAND_111;
  reg  _T_7371; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26962.4]
  reg [31:0] _RAND_112;
  reg  _T_7340; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26920.4]
  reg [31:0] _RAND_113;
  reg  _T_7309; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26878.4]
  reg [31:0] _RAND_114;
  reg  _T_7278; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26836.4]
  reg [31:0] _RAND_115;
  reg  _T_7247; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26794.4]
  reg [31:0] _RAND_116;
  reg  _T_7216; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26752.4]
  reg [31:0] _RAND_117;
  reg  _T_7185; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26710.4]
  reg [31:0] _RAND_118;
  reg  _T_7154; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26668.4]
  reg [31:0] _RAND_119;
  reg  _T_7123; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26626.4]
  reg [31:0] _RAND_120;
  reg  _T_7092; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26584.4]
  reg [31:0] _RAND_121;
  reg  _T_7061; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26542.4]
  reg [31:0] _RAND_122;
  reg  _T_7030; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26500.4]
  reg [31:0] _RAND_123;
  reg  _T_6999; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26458.4]
  reg [31:0] _RAND_124;
  reg  _T_6968; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26416.4]
  reg [31:0] _RAND_125;
  reg  _T_6937; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26374.4]
  reg [31:0] _RAND_126;
  reg  _T_6906; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26332.4]
  reg [31:0] _RAND_127;
  reg  _T_6875; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26290.4]
  reg [31:0] _RAND_128;
  reg  _T_6844; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26248.4]
  reg [31:0] _RAND_129;
  reg  _T_6813; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26206.4]
  reg [31:0] _RAND_130;
  reg  _T_6782; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26164.4]
  reg [31:0] _RAND_131;
  reg  _T_6751; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26122.4]
  reg [31:0] _RAND_132;
  reg  _T_6720; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26080.4]
  reg [31:0] _RAND_133;
  reg  _T_6689; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@26038.4]
  reg [31:0] _RAND_134;
  reg  _T_6658; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25996.4]
  reg [31:0] _RAND_135;
  reg  _T_6627; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25954.4]
  reg [31:0] _RAND_136;
  reg  _T_6596; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25912.4]
  reg [31:0] _RAND_137;
  reg  _T_6565; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25870.4]
  reg [31:0] _RAND_138;
  reg  _T_6534; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25828.4]
  reg [31:0] _RAND_139;
  reg  _T_6503; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25786.4]
  reg [31:0] _RAND_140;
  reg  _T_6472; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25744.4]
  reg [31:0] _RAND_141;
  reg  _T_6441; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25702.4]
  reg [31:0] _RAND_142;
  reg  _T_6410; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25660.4]
  reg [31:0] _RAND_143;
  reg  _T_6379; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25618.4]
  reg [31:0] _RAND_144;
  reg  _T_6348; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25576.4]
  reg [31:0] _RAND_145;
  reg  _T_6317; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25534.4]
  reg [31:0] _RAND_146;
  reg  _T_6286; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25492.4]
  reg [31:0] _RAND_147;
  reg  _T_6255; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25450.4]
  reg [31:0] _RAND_148;
  reg  _T_6224; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25408.4]
  reg [31:0] _RAND_149;
  reg  _T_6193; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25366.4]
  reg [31:0] _RAND_150;
  reg  _T_6162; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25324.4]
  reg [31:0] _RAND_151;
  reg  _T_6131; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25282.4]
  reg [31:0] _RAND_152;
  reg  _T_6100; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25240.4]
  reg [31:0] _RAND_153;
  reg  _T_6069; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25198.4]
  reg [31:0] _RAND_154;
  reg  _T_6038; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25156.4]
  reg [31:0] _RAND_155;
  reg  _T_6007; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25114.4]
  reg [31:0] _RAND_156;
  reg  _T_5976; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25072.4]
  reg [31:0] _RAND_157;
  reg  _T_5945; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@25030.4]
  reg [31:0] _RAND_158;
  reg  _T_5914; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24988.4]
  reg [31:0] _RAND_159;
  reg  _T_5883; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24946.4]
  reg [31:0] _RAND_160;
  reg  _T_5852; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24904.4]
  reg [31:0] _RAND_161;
  reg  _T_5821; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24862.4]
  reg [31:0] _RAND_162;
  reg  _T_5790; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24820.4]
  reg [31:0] _RAND_163;
  reg  _T_5759; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24778.4]
  reg [31:0] _RAND_164;
  reg  _T_5728; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24736.4]
  reg [31:0] _RAND_165;
  reg  _T_5697; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24694.4]
  reg [31:0] _RAND_166;
  reg  _T_5666; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24652.4]
  reg [31:0] _RAND_167;
  reg  _T_5635; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24610.4]
  reg [31:0] _RAND_168;
  reg  _T_5604; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24568.4]
  reg [31:0] _RAND_169;
  reg  _T_5573; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24526.4]
  reg [31:0] _RAND_170;
  reg  _T_5542; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24484.4]
  reg [31:0] _RAND_171;
  reg  _T_5511; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24442.4]
  reg [31:0] _RAND_172;
  reg  _T_5480; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24400.4]
  reg [31:0] _RAND_173;
  reg  _T_5449; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24358.4]
  reg [31:0] _RAND_174;
  reg  _T_5418; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24316.4]
  reg [31:0] _RAND_175;
  reg  _T_5387; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24274.4]
  reg [31:0] _RAND_176;
  reg  _T_5356; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24232.4]
  reg [31:0] _RAND_177;
  reg  _T_5325; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24190.4]
  reg [31:0] _RAND_178;
  reg  _T_5294; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24148.4]
  reg [31:0] _RAND_179;
  reg  _T_5263; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24106.4]
  reg [31:0] _RAND_180;
  reg  _T_5232; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24064.4]
  reg [31:0] _RAND_181;
  reg  _T_5201; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@24022.4]
  reg [31:0] _RAND_182;
  reg  _T_5170; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23980.4]
  reg [31:0] _RAND_183;
  reg  _T_5139; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23938.4]
  reg [31:0] _RAND_184;
  reg  _T_5108; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23896.4]
  reg [31:0] _RAND_185;
  reg  _T_5077; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23854.4]
  reg [31:0] _RAND_186;
  reg  _T_5046; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23812.4]
  reg [31:0] _RAND_187;
  reg  _T_5015; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23770.4]
  reg [31:0] _RAND_188;
  reg  _T_4984; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23728.4]
  reg [31:0] _RAND_189;
  reg  _T_4953; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23686.4]
  reg [31:0] _RAND_190;
  reg  _T_4922; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23644.4]
  reg [31:0] _RAND_191;
  reg  _T_4891; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23602.4]
  reg [31:0] _RAND_192;
  reg  _T_4860; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23560.4]
  reg [31:0] _RAND_193;
  reg  _T_4829; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23518.4]
  reg [31:0] _RAND_194;
  reg  _T_4798; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23476.4]
  reg [31:0] _RAND_195;
  reg  _T_4767; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23434.4]
  reg [31:0] _RAND_196;
  reg  _T_4736; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23392.4]
  reg [31:0] _RAND_197;
  reg  _T_4705; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23350.4]
  reg [31:0] _RAND_198;
  reg  _T_4674; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23308.4]
  reg [31:0] _RAND_199;
  reg  _T_4643; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23266.4]
  reg [31:0] _RAND_200;
  reg  _T_4612; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23224.4]
  reg [31:0] _RAND_201;
  reg  _T_4581; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23182.4]
  reg [31:0] _RAND_202;
  reg  _T_4550; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23140.4]
  reg [31:0] _RAND_203;
  reg  _T_4519; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23098.4]
  reg [31:0] _RAND_204;
  reg  _T_4488; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23056.4]
  reg [31:0] _RAND_205;
  reg  _T_4457; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@23014.4]
  reg [31:0] _RAND_206;
  reg  _T_4426; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22972.4]
  reg [31:0] _RAND_207;
  reg  _T_4395; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22930.4]
  reg [31:0] _RAND_208;
  reg  _T_4364; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22888.4]
  reg [31:0] _RAND_209;
  reg  _T_4333; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22846.4]
  reg [31:0] _RAND_210;
  reg  _T_4302; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22804.4]
  reg [31:0] _RAND_211;
  reg  _T_4271; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22762.4]
  reg [31:0] _RAND_212;
  reg  _T_4240; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22720.4]
  reg [31:0] _RAND_213;
  reg  _T_4209; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22678.4]
  reg [31:0] _RAND_214;
  reg  _T_4178; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22636.4]
  reg [31:0] _RAND_215;
  reg  _T_4147; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22594.4]
  reg [31:0] _RAND_216;
  reg  _T_4116; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22552.4]
  reg [31:0] _RAND_217;
  reg  _T_4085; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22510.4]
  reg [31:0] _RAND_218;
  reg  _T_4054; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22468.4]
  reg [31:0] _RAND_219;
  reg  _T_4023; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22426.4]
  reg [31:0] _RAND_220;
  reg  _T_3992; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22384.4]
  reg [31:0] _RAND_221;
  reg  _T_3961; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22342.4]
  reg [31:0] _RAND_222;
  reg  _T_3930; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22300.4]
  reg [31:0] _RAND_223;
  reg  _T_3899; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22258.4]
  reg [31:0] _RAND_224;
  reg  _T_3868; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22216.4]
  reg [31:0] _RAND_225;
  reg  _T_3837; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22174.4]
  reg [31:0] _RAND_226;
  reg  _T_3806; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22132.4]
  reg [31:0] _RAND_227;
  reg  _T_3775; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22090.4]
  reg [31:0] _RAND_228;
  reg  _T_3744; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22048.4]
  reg [31:0] _RAND_229;
  reg  _T_3713; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@22006.4]
  reg [31:0] _RAND_230;
  reg  _T_3682; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21964.4]
  reg [31:0] _RAND_231;
  reg  _T_3651; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21922.4]
  reg [31:0] _RAND_232;
  reg  _T_3620; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21880.4]
  reg [31:0] _RAND_233;
  reg  _T_3589; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21838.4]
  reg [31:0] _RAND_234;
  reg  _T_3558; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21796.4]
  reg [31:0] _RAND_235;
  reg  _T_3527; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21754.4]
  reg [31:0] _RAND_236;
  reg  _T_3496; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21712.4]
  reg [31:0] _RAND_237;
  reg  _T_3465; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21670.4]
  reg [31:0] _RAND_238;
  reg  _T_3434; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21628.4]
  reg [31:0] _RAND_239;
  reg  _T_3403; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21586.4]
  reg [31:0] _RAND_240;
  reg  _T_3372; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21544.4]
  reg [31:0] _RAND_241;
  reg  _T_3341; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21502.4]
  reg [31:0] _RAND_242;
  reg  _T_3310; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21460.4]
  reg [31:0] _RAND_243;
  reg  _T_3279; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21418.4]
  reg [31:0] _RAND_244;
  reg  _T_3248; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21376.4]
  reg [31:0] _RAND_245;
  reg  _T_3217; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21334.4]
  reg [31:0] _RAND_246;
  reg  _T_3186; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21292.4]
  reg [31:0] _RAND_247;
  reg  _T_3155; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21250.4]
  reg [31:0] _RAND_248;
  reg  _T_3124; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21208.4]
  reg [31:0] _RAND_249;
  reg  _T_3093; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21166.4]
  reg [31:0] _RAND_250;
  reg  _T_3062; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21124.4]
  reg [31:0] _RAND_251;
  reg  _T_3031; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21082.4]
  reg [31:0] _RAND_252;
  reg  _T_3000; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@21040.4]
  reg [31:0] _RAND_253;
  reg  _T_2969; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@20998.4]
  reg [31:0] _RAND_254;
  reg  _T_2938; // @[ToAXI4.scala 225:28:boom.system.TestHarness.MegaBoomConfig.fir@20956.4]
  reg [31:0] _RAND_255;
  wire  _GEN_259; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_260; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_261; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_262; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_263; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_264; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_265; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_266; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_267; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_268; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_269; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_270; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_271; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_272; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_273; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_274; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_275; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_276; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_277; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_278; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_279; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_280; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_281; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_282; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_283; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_284; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_285; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_286; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_287; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_288; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_289; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_290; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_291; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_292; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_293; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_294; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_295; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_296; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_297; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_298; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_299; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_300; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_301; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_302; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_303; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_304; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_305; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_306; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_307; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_308; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_309; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_310; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_311; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_312; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_313; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_314; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_315; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_316; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_317; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_318; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_319; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_320; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_321; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_322; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_323; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_324; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_325; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_326; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_327; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_328; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_329; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_330; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_331; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_332; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_333; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_334; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_335; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_336; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_337; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_338; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_339; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_340; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_341; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_342; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_343; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_344; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_345; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_346; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_347; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_348; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_349; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_350; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_351; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_352; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_353; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_354; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_355; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_356; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_357; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_358; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_359; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_360; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_361; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_362; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_363; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_364; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_365; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_366; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_367; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_368; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_369; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_370; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_371; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_372; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_373; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_374; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_375; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_376; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_377; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_378; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_379; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_380; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_381; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_382; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_383; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_384; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_385; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_386; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_387; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_388; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_389; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_390; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_391; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_392; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_393; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_394; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_395; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_396; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_397; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_398; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_399; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_400; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_401; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_402; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_403; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_404; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_405; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_406; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_407; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_408; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_409; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_410; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_411; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_412; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_413; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_414; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_415; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_416; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_417; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_418; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_419; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_420; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_421; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_422; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_423; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_424; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_425; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_426; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_427; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_428; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_429; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_430; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_431; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_432; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_433; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_434; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_435; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_436; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_437; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_438; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_439; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_440; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_441; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_442; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_443; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_444; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_445; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_446; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_447; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_448; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_449; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_450; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_451; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_452; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_453; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_454; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_455; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_456; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_457; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_458; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_459; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_460; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_461; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_462; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_463; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_464; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_465; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_466; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_467; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_468; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_469; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_470; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_471; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_472; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_473; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_474; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_475; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_476; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_477; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_478; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_479; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_480; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_481; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_482; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_483; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_484; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_485; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_486; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_487; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_488; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_489; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_490; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_491; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_492; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_493; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_494; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_495; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_496; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_497; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_498; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_499; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_500; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_501; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_502; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_503; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_504; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_505; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_506; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_507; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_508; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_509; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_510; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_511; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_512; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _GEN_513; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  reg [2:0] _T_2307; // @[Edges.scala 229:27:boom.system.TestHarness.MegaBoomConfig.fir@20243.4]
  reg [31:0] _RAND_256;
  wire  _T_2311; // @[Edges.scala 231:25:boom.system.TestHarness.MegaBoomConfig.fir@20247.4]
  wire  _T_2377; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  wire  _T_2378; // @[ToAXI4.scala 177:21:boom.system.TestHarness.MegaBoomConfig.fir@20364.4]
  reg  _T_2365; // @[ToAXI4.scala 160:30:boom.system.TestHarness.MegaBoomConfig.fir@20339.4]
  reg [31:0] _RAND_257;
  wire  _T_2338_ready; // @[ToAXI4.scala 146:25:boom.system.TestHarness.MegaBoomConfig.fir@20281.4 Decoupled.scala 296:17:boom.system.TestHarness.MegaBoomConfig.fir@20315.4]
  wire  _T_2379; // @[ToAXI4.scala 177:52:boom.system.TestHarness.MegaBoomConfig.fir@20365.4]
  wire  _T_2341_ready; // @[ToAXI4.scala 147:23:boom.system.TestHarness.MegaBoomConfig.fir@20283.4 Decoupled.scala 296:17:boom.system.TestHarness.MegaBoomConfig.fir@20292.4]
  wire  _T_2380; // @[ToAXI4.scala 177:70:boom.system.TestHarness.MegaBoomConfig.fir@20366.4]
  wire  _T_2381; // @[ToAXI4.scala 177:34:boom.system.TestHarness.MegaBoomConfig.fir@20367.4]
  wire  _T_2382; // @[ToAXI4.scala 177:28:boom.system.TestHarness.MegaBoomConfig.fir@20368.4]
  wire  _T_2297; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@20234.4]
  wire [12:0] _T_2299; // @[package.scala 185:77:boom.system.TestHarness.MegaBoomConfig.fir@20236.4]
  wire [5:0] _T_2300; // @[package.scala 185:82:boom.system.TestHarness.MegaBoomConfig.fir@20237.4]
  wire [5:0] _T_2301; // @[package.scala 185:46:boom.system.TestHarness.MegaBoomConfig.fir@20238.4]
  wire [2:0] _T_2302; // @[Edges.scala 220:59:boom.system.TestHarness.MegaBoomConfig.fir@20239.4]
  wire [2:0] _T_2305; // @[Edges.scala 221:14:boom.system.TestHarness.MegaBoomConfig.fir@20242.4]
  wire [3:0] _T_2308; // @[Edges.scala 230:28:boom.system.TestHarness.MegaBoomConfig.fir@20244.4]
  wire [3:0] _T_2309; // @[Edges.scala 230:28:boom.system.TestHarness.MegaBoomConfig.fir@20245.4]
  wire [2:0] _T_2310; // @[Edges.scala 230:28:boom.system.TestHarness.MegaBoomConfig.fir@20246.4]
  wire  _T_2312; // @[Edges.scala 232:25:boom.system.TestHarness.MegaBoomConfig.fir@20248.4]
  wire  _T_2313; // @[Edges.scala 232:47:boom.system.TestHarness.MegaBoomConfig.fir@20249.4]
  wire  _T_2314; // @[Edges.scala 232:37:boom.system.TestHarness.MegaBoomConfig.fir@20250.4]
  wire [10:0] _GEN_773; // @[ToAXI4.scala 134:55:boom.system.TestHarness.MegaBoomConfig.fir@20275.4]
  wire [10:0] _T_2328; // @[ToAXI4.scala 134:55:boom.system.TestHarness.MegaBoomConfig.fir@20275.4]
  wire [10:0] _GEN_774; // @[ToAXI4.scala 134:45:boom.system.TestHarness.MegaBoomConfig.fir@20276.4]
  wire [10:0] _T_2329; // @[ToAXI4.scala 134:45:boom.system.TestHarness.MegaBoomConfig.fir@20276.4]
  wire [7:0] _T_2330; // @[ToAXI4.scala 137:50:boom.system.TestHarness.MegaBoomConfig.fir@20277.4]
  wire [2:0] _T_2331; // @[ToAXI4.scala 138:50:boom.system.TestHarness.MegaBoomConfig.fir@20278.4]
  wire [7:0] _T_2332; // @[ToAXI4.scala 141:50:boom.system.TestHarness.MegaBoomConfig.fir@20279.4]
  wire [2:0] _T_2333; // @[ToAXI4.scala 142:50:boom.system.TestHarness.MegaBoomConfig.fir@20280.4]
  wire  _T_2356_bits_wen; // @[Decoupled.scala 314:19:boom.system.TestHarness.MegaBoomConfig.fir@20316.4 Decoupled.scala 315:14:boom.system.TestHarness.MegaBoomConfig.fir@20317.4]
  wire  _T_2360; // @[ToAXI4.scala 154:42:boom.system.TestHarness.MegaBoomConfig.fir@20332.4]
  wire  _T_2356_valid; // @[Decoupled.scala 314:19:boom.system.TestHarness.MegaBoomConfig.fir@20316.4 Decoupled.scala 316:15:boom.system.TestHarness.MegaBoomConfig.fir@20328.4]
  wire  _T_2367; // @[ToAXI4.scala 161:38:boom.system.TestHarness.MegaBoomConfig.fir@20342.6]
  wire [7:0] _GEN_3; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_4; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_5; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_6; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_7; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_8; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_9; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_10; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_11; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_12; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_13; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_14; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_15; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_16; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_17; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_18; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_19; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_20; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_21; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_22; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_23; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_24; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_25; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_26; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_27; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_28; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_29; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_30; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_31; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_32; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_33; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_34; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_35; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_36; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_37; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_38; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_39; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_40; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_41; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_42; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_43; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_44; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_45; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_46; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_47; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_48; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_49; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_50; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_51; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_52; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_53; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_54; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_55; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_56; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_57; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_58; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_59; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_60; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_61; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_62; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_63; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_64; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_65; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_66; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_67; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_68; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_69; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_70; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_71; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_72; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_73; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_74; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_75; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_76; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_77; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_78; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_79; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_80; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_81; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_82; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_83; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_84; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_85; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_86; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_87; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_88; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_89; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_90; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_91; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_92; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_93; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_94; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_95; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_96; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_97; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_98; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_99; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_100; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_101; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_102; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_103; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_104; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_105; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_106; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_107; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_108; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_109; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_110; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_111; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_112; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_113; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_114; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_115; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_116; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_117; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_118; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_119; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_120; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_121; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_122; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_123; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_124; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_125; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_126; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_127; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_128; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_129; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_130; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_131; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_132; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_133; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_134; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_135; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_136; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_137; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_138; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_139; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_140; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_141; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_142; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_143; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_144; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_145; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_146; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_147; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_148; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_149; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_150; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_151; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_152; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_153; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_154; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_155; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_156; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_157; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_158; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_159; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_160; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_161; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_162; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_163; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_164; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_165; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_166; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_167; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_168; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_169; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_170; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_171; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_172; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_173; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_174; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_175; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_176; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_177; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_178; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_179; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_180; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_181; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_182; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_183; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_184; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_185; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_186; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_187; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_188; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_189; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_190; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_191; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_192; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_193; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_194; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_195; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_196; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_197; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_198; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_199; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_200; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_201; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_202; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_203; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_204; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_205; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_206; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_207; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_208; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_209; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_210; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_211; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_212; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_213; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_214; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_215; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_216; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_217; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_218; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_219; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_220; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_221; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_222; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_223; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_224; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_225; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_226; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_227; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_228; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_229; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_230; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_231; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_232; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_233; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_234; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_235; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_236; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_237; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_238; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_239; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_240; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_241; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_242; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_243; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_244; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_245; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_246; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_247; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_248; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_249; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_250; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_251; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_252; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_253; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_254; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_255; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_256; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [7:0] _GEN_257; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  wire [17:0] _T_2370; // @[package.scala 185:77:boom.system.TestHarness.MegaBoomConfig.fir@20349.4]
  wire [10:0] _T_2371; // @[package.scala 185:82:boom.system.TestHarness.MegaBoomConfig.fir@20350.4]
  wire [10:0] _T_2372; // @[package.scala 185:46:boom.system.TestHarness.MegaBoomConfig.fir@20351.4]
  wire  _T_2374; // @[ToAXI4.scala 168:31:boom.system.TestHarness.MegaBoomConfig.fir@20354.4]
  wire  _T_2384; // @[ToAXI4.scala 178:31:boom.system.TestHarness.MegaBoomConfig.fir@20371.4]
  wire  _T_2385; // @[ToAXI4.scala 178:61:boom.system.TestHarness.MegaBoomConfig.fir@20372.4]
  wire  _T_2386; // @[ToAXI4.scala 178:69:boom.system.TestHarness.MegaBoomConfig.fir@20373.4]
  wire  _T_2387; // @[ToAXI4.scala 178:51:boom.system.TestHarness.MegaBoomConfig.fir@20374.4]
  wire  _T_2388; // @[ToAXI4.scala 178:45:boom.system.TestHarness.MegaBoomConfig.fir@20375.4]
  wire  _T_2391; // @[ToAXI4.scala 180:43:boom.system.TestHarness.MegaBoomConfig.fir@20379.4]
  reg  _T_2395; // @[ToAXI4.scala 187:30:boom.system.TestHarness.MegaBoomConfig.fir@20386.4]
  reg [31:0] _RAND_258;
  wire  _T_2396; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@20387.4]
  wire  _T_2397; // @[ToAXI4.scala 188:42:boom.system.TestHarness.MegaBoomConfig.fir@20389.6]
  wire  _T_2398; // @[ToAXI4.scala 190:32:boom.system.TestHarness.MegaBoomConfig.fir@20392.4]
  wire  _T_2399; // @[ToAXI4.scala 193:36:boom.system.TestHarness.MegaBoomConfig.fir@20394.4]
  wire  _T_2401; // @[ToAXI4.scala 194:24:boom.system.TestHarness.MegaBoomConfig.fir@20397.4]
  reg  _T_2403; // @[ToAXI4.scala 199:28:boom.system.TestHarness.MegaBoomConfig.fir@20399.4]
  reg [31:0] _RAND_259;
  wire  _T_2405; // @[ToAXI4.scala 201:39:boom.system.TestHarness.MegaBoomConfig.fir@20404.4]
  reg  _T_2407; // @[Reg.scala 11:16:boom.system.TestHarness.MegaBoomConfig.fir@20405.4]
  reg [31:0] _RAND_260;
  wire  _GEN_516; // @[Reg.scala 12:19:boom.system.TestHarness.MegaBoomConfig.fir@20406.4]
  wire  _T_2409; // @[ToAXI4.scala 202:39:boom.system.TestHarness.MegaBoomConfig.fir@20410.4]
  wire  _T_2410; // @[ToAXI4.scala 203:39:boom.system.TestHarness.MegaBoomConfig.fir@20411.4]
  wire  _T_2411; // @[ToAXI4.scala 205:100:boom.system.TestHarness.MegaBoomConfig.fir@20412.4]
  wire [255:0] _T_2418; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@20437.4]
  wire  _T_2420; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20439.4]
  wire  _T_2421; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20440.4]
  wire  _T_2422; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20441.4]
  wire  _T_2423; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20442.4]
  wire  _T_2424; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20443.4]
  wire  _T_2425; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20444.4]
  wire  _T_2426; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20445.4]
  wire  _T_2427; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20446.4]
  wire  _T_2428; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20447.4]
  wire  _T_2429; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20448.4]
  wire  _T_2430; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20449.4]
  wire  _T_2431; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20450.4]
  wire  _T_2432; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20451.4]
  wire  _T_2433; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20452.4]
  wire  _T_2434; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20453.4]
  wire  _T_2435; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20454.4]
  wire  _T_2436; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20455.4]
  wire  _T_2437; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20456.4]
  wire  _T_2438; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20457.4]
  wire  _T_2439; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20458.4]
  wire  _T_2440; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20459.4]
  wire  _T_2441; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20460.4]
  wire  _T_2442; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20461.4]
  wire  _T_2443; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20462.4]
  wire  _T_2444; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20463.4]
  wire  _T_2445; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20464.4]
  wire  _T_2446; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20465.4]
  wire  _T_2447; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20466.4]
  wire  _T_2448; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20467.4]
  wire  _T_2449; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20468.4]
  wire  _T_2450; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20469.4]
  wire  _T_2451; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20470.4]
  wire  _T_2452; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20471.4]
  wire  _T_2453; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20472.4]
  wire  _T_2454; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20473.4]
  wire  _T_2455; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20474.4]
  wire  _T_2456; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20475.4]
  wire  _T_2457; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20476.4]
  wire  _T_2458; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20477.4]
  wire  _T_2459; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20478.4]
  wire  _T_2460; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20479.4]
  wire  _T_2461; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20480.4]
  wire  _T_2462; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20481.4]
  wire  _T_2463; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20482.4]
  wire  _T_2464; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20483.4]
  wire  _T_2465; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20484.4]
  wire  _T_2466; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20485.4]
  wire  _T_2467; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20486.4]
  wire  _T_2468; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20487.4]
  wire  _T_2469; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20488.4]
  wire  _T_2470; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20489.4]
  wire  _T_2471; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20490.4]
  wire  _T_2472; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20491.4]
  wire  _T_2473; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20492.4]
  wire  _T_2474; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20493.4]
  wire  _T_2475; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20494.4]
  wire  _T_2476; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20495.4]
  wire  _T_2477; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20496.4]
  wire  _T_2478; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20497.4]
  wire  _T_2479; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20498.4]
  wire  _T_2480; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20499.4]
  wire  _T_2481; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20500.4]
  wire  _T_2482; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20501.4]
  wire  _T_2483; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20502.4]
  wire  _T_2484; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20503.4]
  wire  _T_2485; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20504.4]
  wire  _T_2486; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20505.4]
  wire  _T_2487; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20506.4]
  wire  _T_2488; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20507.4]
  wire  _T_2489; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20508.4]
  wire  _T_2490; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20509.4]
  wire  _T_2491; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20510.4]
  wire  _T_2492; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20511.4]
  wire  _T_2493; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20512.4]
  wire  _T_2494; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20513.4]
  wire  _T_2495; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20514.4]
  wire  _T_2496; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20515.4]
  wire  _T_2497; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20516.4]
  wire  _T_2498; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20517.4]
  wire  _T_2499; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20518.4]
  wire  _T_2500; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20519.4]
  wire  _T_2501; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20520.4]
  wire  _T_2502; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20521.4]
  wire  _T_2503; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20522.4]
  wire  _T_2504; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20523.4]
  wire  _T_2505; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20524.4]
  wire  _T_2506; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20525.4]
  wire  _T_2507; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20526.4]
  wire  _T_2508; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20527.4]
  wire  _T_2509; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20528.4]
  wire  _T_2510; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20529.4]
  wire  _T_2511; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20530.4]
  wire  _T_2512; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20531.4]
  wire  _T_2513; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20532.4]
  wire  _T_2514; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20533.4]
  wire  _T_2515; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20534.4]
  wire  _T_2516; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20535.4]
  wire  _T_2517; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20536.4]
  wire  _T_2518; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20537.4]
  wire  _T_2519; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20538.4]
  wire  _T_2520; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20539.4]
  wire  _T_2521; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20540.4]
  wire  _T_2522; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20541.4]
  wire  _T_2523; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20542.4]
  wire  _T_2524; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20543.4]
  wire  _T_2525; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20544.4]
  wire  _T_2526; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20545.4]
  wire  _T_2527; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20546.4]
  wire  _T_2528; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20547.4]
  wire  _T_2529; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20548.4]
  wire  _T_2530; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20549.4]
  wire  _T_2531; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20550.4]
  wire  _T_2532; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20551.4]
  wire  _T_2533; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20552.4]
  wire  _T_2534; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20553.4]
  wire  _T_2535; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20554.4]
  wire  _T_2536; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20555.4]
  wire  _T_2537; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20556.4]
  wire  _T_2538; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20557.4]
  wire  _T_2539; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20558.4]
  wire  _T_2540; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20559.4]
  wire  _T_2541; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20560.4]
  wire  _T_2542; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20561.4]
  wire  _T_2543; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20562.4]
  wire  _T_2544; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20563.4]
  wire  _T_2545; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20564.4]
  wire  _T_2546; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20565.4]
  wire  _T_2547; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20566.4]
  wire  _T_2548; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20567.4]
  wire  _T_2549; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20568.4]
  wire  _T_2550; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20569.4]
  wire  _T_2551; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20570.4]
  wire  _T_2552; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20571.4]
  wire  _T_2553; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20572.4]
  wire  _T_2554; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20573.4]
  wire  _T_2555; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20574.4]
  wire  _T_2556; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20575.4]
  wire  _T_2557; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20576.4]
  wire  _T_2558; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20577.4]
  wire  _T_2559; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20578.4]
  wire  _T_2560; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20579.4]
  wire  _T_2561; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20580.4]
  wire  _T_2562; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20581.4]
  wire  _T_2563; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20582.4]
  wire  _T_2564; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20583.4]
  wire  _T_2565; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20584.4]
  wire  _T_2566; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20585.4]
  wire  _T_2567; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20586.4]
  wire  _T_2568; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20587.4]
  wire  _T_2569; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20588.4]
  wire  _T_2570; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20589.4]
  wire  _T_2571; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20590.4]
  wire  _T_2572; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20591.4]
  wire  _T_2573; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20592.4]
  wire  _T_2574; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20593.4]
  wire  _T_2575; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20594.4]
  wire  _T_2576; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20595.4]
  wire  _T_2577; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20596.4]
  wire  _T_2578; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20597.4]
  wire  _T_2579; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20598.4]
  wire  _T_2580; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20599.4]
  wire  _T_2581; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20600.4]
  wire  _T_2582; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20601.4]
  wire  _T_2583; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20602.4]
  wire  _T_2584; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20603.4]
  wire  _T_2585; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20604.4]
  wire  _T_2586; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20605.4]
  wire  _T_2587; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20606.4]
  wire  _T_2588; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20607.4]
  wire  _T_2589; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20608.4]
  wire  _T_2590; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20609.4]
  wire  _T_2591; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20610.4]
  wire  _T_2592; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20611.4]
  wire  _T_2593; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20612.4]
  wire  _T_2594; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20613.4]
  wire  _T_2595; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20614.4]
  wire  _T_2596; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20615.4]
  wire  _T_2597; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20616.4]
  wire  _T_2598; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20617.4]
  wire  _T_2599; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20618.4]
  wire  _T_2600; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20619.4]
  wire  _T_2601; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20620.4]
  wire  _T_2602; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20621.4]
  wire  _T_2603; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20622.4]
  wire  _T_2604; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20623.4]
  wire  _T_2605; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20624.4]
  wire  _T_2606; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20625.4]
  wire  _T_2607; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20626.4]
  wire  _T_2608; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20627.4]
  wire  _T_2609; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20628.4]
  wire  _T_2610; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20629.4]
  wire  _T_2611; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20630.4]
  wire  _T_2612; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20631.4]
  wire  _T_2613; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20632.4]
  wire  _T_2614; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20633.4]
  wire  _T_2615; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20634.4]
  wire  _T_2616; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20635.4]
  wire  _T_2617; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20636.4]
  wire  _T_2618; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20637.4]
  wire  _T_2619; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20638.4]
  wire  _T_2620; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20639.4]
  wire  _T_2621; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20640.4]
  wire  _T_2622; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20641.4]
  wire  _T_2623; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20642.4]
  wire  _T_2624; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20643.4]
  wire  _T_2625; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20644.4]
  wire  _T_2626; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20645.4]
  wire  _T_2627; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20646.4]
  wire  _T_2628; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20647.4]
  wire  _T_2629; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20648.4]
  wire  _T_2630; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20649.4]
  wire  _T_2631; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20650.4]
  wire  _T_2632; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20651.4]
  wire  _T_2633; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20652.4]
  wire  _T_2634; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20653.4]
  wire  _T_2635; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20654.4]
  wire  _T_2636; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20655.4]
  wire  _T_2637; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20656.4]
  wire  _T_2638; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20657.4]
  wire  _T_2639; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20658.4]
  wire  _T_2640; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20659.4]
  wire  _T_2641; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20660.4]
  wire  _T_2642; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20661.4]
  wire  _T_2643; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20662.4]
  wire  _T_2644; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20663.4]
  wire  _T_2645; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20664.4]
  wire  _T_2646; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20665.4]
  wire  _T_2647; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20666.4]
  wire  _T_2648; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20667.4]
  wire  _T_2649; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20668.4]
  wire  _T_2650; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20669.4]
  wire  _T_2651; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20670.4]
  wire  _T_2652; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20671.4]
  wire  _T_2653; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20672.4]
  wire  _T_2654; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20673.4]
  wire  _T_2655; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20674.4]
  wire  _T_2656; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20675.4]
  wire  _T_2657; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20676.4]
  wire  _T_2658; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20677.4]
  wire  _T_2659; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20678.4]
  wire  _T_2660; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20679.4]
  wire  _T_2661; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20680.4]
  wire  _T_2662; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20681.4]
  wire  _T_2663; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20682.4]
  wire  _T_2664; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20683.4]
  wire  _T_2665; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20684.4]
  wire  _T_2666; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20685.4]
  wire  _T_2667; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20686.4]
  wire  _T_2668; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20687.4]
  wire  _T_2669; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20688.4]
  wire  _T_2670; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20689.4]
  wire  _T_2671; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20690.4]
  wire  _T_2672; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20691.4]
  wire  _T_2673; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20692.4]
  wire  _T_2674; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20693.4]
  wire  _T_2675; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20694.4]
  wire [7:0] _T_2676; // @[ToAXI4.scala 214:31:boom.system.TestHarness.MegaBoomConfig.fir@20695.4]
  wire [255:0] _T_2678; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@20697.4]
  wire  _T_2680; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20699.4]
  wire  _T_2681; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20700.4]
  wire  _T_2682; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20701.4]
  wire  _T_2683; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20702.4]
  wire  _T_2684; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20703.4]
  wire  _T_2685; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20704.4]
  wire  _T_2686; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20705.4]
  wire  _T_2687; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20706.4]
  wire  _T_2688; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20707.4]
  wire  _T_2689; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20708.4]
  wire  _T_2690; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20709.4]
  wire  _T_2691; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20710.4]
  wire  _T_2692; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20711.4]
  wire  _T_2693; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20712.4]
  wire  _T_2694; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20713.4]
  wire  _T_2695; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20714.4]
  wire  _T_2696; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20715.4]
  wire  _T_2697; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20716.4]
  wire  _T_2698; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20717.4]
  wire  _T_2699; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20718.4]
  wire  _T_2700; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20719.4]
  wire  _T_2701; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20720.4]
  wire  _T_2702; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20721.4]
  wire  _T_2703; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20722.4]
  wire  _T_2704; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20723.4]
  wire  _T_2705; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20724.4]
  wire  _T_2706; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20725.4]
  wire  _T_2707; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20726.4]
  wire  _T_2708; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20727.4]
  wire  _T_2709; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20728.4]
  wire  _T_2710; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20729.4]
  wire  _T_2711; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20730.4]
  wire  _T_2712; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20731.4]
  wire  _T_2713; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20732.4]
  wire  _T_2714; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20733.4]
  wire  _T_2715; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20734.4]
  wire  _T_2716; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20735.4]
  wire  _T_2717; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20736.4]
  wire  _T_2718; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20737.4]
  wire  _T_2719; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20738.4]
  wire  _T_2720; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20739.4]
  wire  _T_2721; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20740.4]
  wire  _T_2722; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20741.4]
  wire  _T_2723; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20742.4]
  wire  _T_2724; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20743.4]
  wire  _T_2725; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20744.4]
  wire  _T_2726; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20745.4]
  wire  _T_2727; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20746.4]
  wire  _T_2728; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20747.4]
  wire  _T_2729; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20748.4]
  wire  _T_2730; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20749.4]
  wire  _T_2731; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20750.4]
  wire  _T_2732; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20751.4]
  wire  _T_2733; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20752.4]
  wire  _T_2734; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20753.4]
  wire  _T_2735; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20754.4]
  wire  _T_2736; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20755.4]
  wire  _T_2737; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20756.4]
  wire  _T_2738; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20757.4]
  wire  _T_2739; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20758.4]
  wire  _T_2740; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20759.4]
  wire  _T_2741; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20760.4]
  wire  _T_2742; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20761.4]
  wire  _T_2743; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20762.4]
  wire  _T_2744; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20763.4]
  wire  _T_2745; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20764.4]
  wire  _T_2746; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20765.4]
  wire  _T_2747; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20766.4]
  wire  _T_2748; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20767.4]
  wire  _T_2749; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20768.4]
  wire  _T_2750; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20769.4]
  wire  _T_2751; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20770.4]
  wire  _T_2752; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20771.4]
  wire  _T_2753; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20772.4]
  wire  _T_2754; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20773.4]
  wire  _T_2755; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20774.4]
  wire  _T_2756; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20775.4]
  wire  _T_2757; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20776.4]
  wire  _T_2758; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20777.4]
  wire  _T_2759; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20778.4]
  wire  _T_2760; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20779.4]
  wire  _T_2761; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20780.4]
  wire  _T_2762; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20781.4]
  wire  _T_2763; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20782.4]
  wire  _T_2764; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20783.4]
  wire  _T_2765; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20784.4]
  wire  _T_2766; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20785.4]
  wire  _T_2767; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20786.4]
  wire  _T_2768; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20787.4]
  wire  _T_2769; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20788.4]
  wire  _T_2770; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20789.4]
  wire  _T_2771; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20790.4]
  wire  _T_2772; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20791.4]
  wire  _T_2773; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20792.4]
  wire  _T_2774; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20793.4]
  wire  _T_2775; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20794.4]
  wire  _T_2776; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20795.4]
  wire  _T_2777; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20796.4]
  wire  _T_2778; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20797.4]
  wire  _T_2779; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20798.4]
  wire  _T_2780; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20799.4]
  wire  _T_2781; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20800.4]
  wire  _T_2782; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20801.4]
  wire  _T_2783; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20802.4]
  wire  _T_2784; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20803.4]
  wire  _T_2785; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20804.4]
  wire  _T_2786; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20805.4]
  wire  _T_2787; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20806.4]
  wire  _T_2788; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20807.4]
  wire  _T_2789; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20808.4]
  wire  _T_2790; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20809.4]
  wire  _T_2791; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20810.4]
  wire  _T_2792; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20811.4]
  wire  _T_2793; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20812.4]
  wire  _T_2794; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20813.4]
  wire  _T_2795; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20814.4]
  wire  _T_2796; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20815.4]
  wire  _T_2797; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20816.4]
  wire  _T_2798; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20817.4]
  wire  _T_2799; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20818.4]
  wire  _T_2800; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20819.4]
  wire  _T_2801; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20820.4]
  wire  _T_2802; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20821.4]
  wire  _T_2803; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20822.4]
  wire  _T_2804; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20823.4]
  wire  _T_2805; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20824.4]
  wire  _T_2806; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20825.4]
  wire  _T_2807; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20826.4]
  wire  _T_2808; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20827.4]
  wire  _T_2809; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20828.4]
  wire  _T_2810; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20829.4]
  wire  _T_2811; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20830.4]
  wire  _T_2812; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20831.4]
  wire  _T_2813; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20832.4]
  wire  _T_2814; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20833.4]
  wire  _T_2815; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20834.4]
  wire  _T_2816; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20835.4]
  wire  _T_2817; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20836.4]
  wire  _T_2818; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20837.4]
  wire  _T_2819; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20838.4]
  wire  _T_2820; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20839.4]
  wire  _T_2821; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20840.4]
  wire  _T_2822; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20841.4]
  wire  _T_2823; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20842.4]
  wire  _T_2824; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20843.4]
  wire  _T_2825; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20844.4]
  wire  _T_2826; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20845.4]
  wire  _T_2827; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20846.4]
  wire  _T_2828; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20847.4]
  wire  _T_2829; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20848.4]
  wire  _T_2830; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20849.4]
  wire  _T_2831; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20850.4]
  wire  _T_2832; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20851.4]
  wire  _T_2833; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20852.4]
  wire  _T_2834; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20853.4]
  wire  _T_2835; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20854.4]
  wire  _T_2836; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20855.4]
  wire  _T_2837; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20856.4]
  wire  _T_2838; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20857.4]
  wire  _T_2839; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20858.4]
  wire  _T_2840; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20859.4]
  wire  _T_2841; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20860.4]
  wire  _T_2842; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20861.4]
  wire  _T_2843; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20862.4]
  wire  _T_2844; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20863.4]
  wire  _T_2845; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20864.4]
  wire  _T_2846; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20865.4]
  wire  _T_2847; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20866.4]
  wire  _T_2848; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20867.4]
  wire  _T_2849; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20868.4]
  wire  _T_2850; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20869.4]
  wire  _T_2851; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20870.4]
  wire  _T_2852; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20871.4]
  wire  _T_2853; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20872.4]
  wire  _T_2854; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20873.4]
  wire  _T_2855; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20874.4]
  wire  _T_2856; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20875.4]
  wire  _T_2857; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20876.4]
  wire  _T_2858; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20877.4]
  wire  _T_2859; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20878.4]
  wire  _T_2860; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20879.4]
  wire  _T_2861; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20880.4]
  wire  _T_2862; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20881.4]
  wire  _T_2863; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20882.4]
  wire  _T_2864; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20883.4]
  wire  _T_2865; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20884.4]
  wire  _T_2866; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20885.4]
  wire  _T_2867; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20886.4]
  wire  _T_2868; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20887.4]
  wire  _T_2869; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20888.4]
  wire  _T_2870; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20889.4]
  wire  _T_2871; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20890.4]
  wire  _T_2872; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20891.4]
  wire  _T_2873; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20892.4]
  wire  _T_2874; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20893.4]
  wire  _T_2875; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20894.4]
  wire  _T_2876; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20895.4]
  wire  _T_2877; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20896.4]
  wire  _T_2878; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20897.4]
  wire  _T_2879; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20898.4]
  wire  _T_2880; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20899.4]
  wire  _T_2881; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20900.4]
  wire  _T_2882; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20901.4]
  wire  _T_2883; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20902.4]
  wire  _T_2884; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20903.4]
  wire  _T_2885; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20904.4]
  wire  _T_2886; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20905.4]
  wire  _T_2887; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20906.4]
  wire  _T_2888; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20907.4]
  wire  _T_2889; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20908.4]
  wire  _T_2890; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20909.4]
  wire  _T_2891; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20910.4]
  wire  _T_2892; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20911.4]
  wire  _T_2893; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20912.4]
  wire  _T_2894; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20913.4]
  wire  _T_2895; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20914.4]
  wire  _T_2896; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20915.4]
  wire  _T_2897; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20916.4]
  wire  _T_2898; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20917.4]
  wire  _T_2899; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20918.4]
  wire  _T_2900; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20919.4]
  wire  _T_2901; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20920.4]
  wire  _T_2902; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20921.4]
  wire  _T_2903; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20922.4]
  wire  _T_2904; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20923.4]
  wire  _T_2905; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20924.4]
  wire  _T_2906; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20925.4]
  wire  _T_2907; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20926.4]
  wire  _T_2908; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20927.4]
  wire  _T_2909; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20928.4]
  wire  _T_2910; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20929.4]
  wire  _T_2911; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20930.4]
  wire  _T_2912; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20931.4]
  wire  _T_2913; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20932.4]
  wire  _T_2914; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20933.4]
  wire  _T_2915; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20934.4]
  wire  _T_2916; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20935.4]
  wire  _T_2917; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20936.4]
  wire  _T_2918; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20937.4]
  wire  _T_2919; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20938.4]
  wire  _T_2920; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20939.4]
  wire  _T_2921; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20940.4]
  wire  _T_2922; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20941.4]
  wire  _T_2923; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20942.4]
  wire  _T_2924; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20943.4]
  wire  _T_2925; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20944.4]
  wire  _T_2926; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20945.4]
  wire  _T_2927; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20946.4]
  wire  _T_2928; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20947.4]
  wire  _T_2929; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20948.4]
  wire  _T_2930; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20949.4]
  wire  _T_2931; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20950.4]
  wire  _T_2932; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20951.4]
  wire  _T_2933; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20952.4]
  wire  _T_2934; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20953.4]
  wire  _T_2935; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20954.4]
  wire  _T_2936; // @[ToAXI4.scala 215:23:boom.system.TestHarness.MegaBoomConfig.fir@20955.4]
  wire  _T_2942; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@20959.4]
  wire  _T_2943; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@20960.4]
  wire  _T_2944; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@20961.4]
  wire  _T_2945; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@20962.4]
  wire  _T_2946; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@20963.4]
  wire  _T_2948; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@20965.4]
  wire [1:0] _T_2949; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@20966.4]
  wire [1:0] _T_2950; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@20967.4]
  wire  _T_2951; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@20968.4]
  wire  _T_2952; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@20970.4]
  wire  _T_2954; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@20972.4]
  wire  _T_2956; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@20974.4]
  wire  _T_2957; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@20975.4]
  wire  _T_2958; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@20980.4]
  wire  _T_2959; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@20981.4]
  wire  _T_2960; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@20982.4]
  wire  _T_2962; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@20984.4]
  wire  _T_2963; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@20985.4]
  wire  _T_2974; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21002.4]
  wire  _T_2975; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21003.4]
  wire  _T_2977; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21005.4]
  wire  _T_2979; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21007.4]
  wire [1:0] _T_2980; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21008.4]
  wire [1:0] _T_2981; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21009.4]
  wire  _T_2982; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21010.4]
  wire  _T_2983; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21012.4]
  wire  _T_2985; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21014.4]
  wire  _T_2987; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21016.4]
  wire  _T_2988; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21017.4]
  wire  _T_2989; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21022.4]
  wire  _T_2990; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21023.4]
  wire  _T_2991; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21024.4]
  wire  _T_2993; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21026.4]
  wire  _T_2994; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21027.4]
  wire  _T_3005; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21044.4]
  wire  _T_3006; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21045.4]
  wire  _T_3008; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21047.4]
  wire  _T_3010; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21049.4]
  wire [1:0] _T_3011; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21050.4]
  wire [1:0] _T_3012; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21051.4]
  wire  _T_3013; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21052.4]
  wire  _T_3014; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21054.4]
  wire  _T_3016; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21056.4]
  wire  _T_3018; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21058.4]
  wire  _T_3019; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21059.4]
  wire  _T_3020; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21064.4]
  wire  _T_3021; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21065.4]
  wire  _T_3022; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21066.4]
  wire  _T_3024; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21068.4]
  wire  _T_3025; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21069.4]
  wire  _T_3036; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21086.4]
  wire  _T_3037; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21087.4]
  wire  _T_3039; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21089.4]
  wire  _T_3041; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21091.4]
  wire [1:0] _T_3042; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21092.4]
  wire [1:0] _T_3043; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21093.4]
  wire  _T_3044; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21094.4]
  wire  _T_3045; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21096.4]
  wire  _T_3047; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21098.4]
  wire  _T_3049; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21100.4]
  wire  _T_3050; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21101.4]
  wire  _T_3051; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21106.4]
  wire  _T_3052; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21107.4]
  wire  _T_3053; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21108.4]
  wire  _T_3055; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21110.4]
  wire  _T_3056; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21111.4]
  wire  _T_3067; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21128.4]
  wire  _T_3068; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21129.4]
  wire  _T_3070; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21131.4]
  wire  _T_3072; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21133.4]
  wire [1:0] _T_3073; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21134.4]
  wire [1:0] _T_3074; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21135.4]
  wire  _T_3075; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21136.4]
  wire  _T_3076; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21138.4]
  wire  _T_3078; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21140.4]
  wire  _T_3080; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21142.4]
  wire  _T_3081; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21143.4]
  wire  _T_3082; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21148.4]
  wire  _T_3083; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21149.4]
  wire  _T_3084; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21150.4]
  wire  _T_3086; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21152.4]
  wire  _T_3087; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21153.4]
  wire  _T_3098; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21170.4]
  wire  _T_3099; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21171.4]
  wire  _T_3101; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21173.4]
  wire  _T_3103; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21175.4]
  wire [1:0] _T_3104; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21176.4]
  wire [1:0] _T_3105; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21177.4]
  wire  _T_3106; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21178.4]
  wire  _T_3107; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21180.4]
  wire  _T_3109; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21182.4]
  wire  _T_3111; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21184.4]
  wire  _T_3112; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21185.4]
  wire  _T_3113; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21190.4]
  wire  _T_3114; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21191.4]
  wire  _T_3115; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21192.4]
  wire  _T_3117; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21194.4]
  wire  _T_3118; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21195.4]
  wire  _T_3129; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21212.4]
  wire  _T_3130; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21213.4]
  wire  _T_3132; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21215.4]
  wire  _T_3134; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21217.4]
  wire [1:0] _T_3135; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21218.4]
  wire [1:0] _T_3136; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21219.4]
  wire  _T_3137; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21220.4]
  wire  _T_3138; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21222.4]
  wire  _T_3140; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21224.4]
  wire  _T_3142; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21226.4]
  wire  _T_3143; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21227.4]
  wire  _T_3144; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21232.4]
  wire  _T_3145; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21233.4]
  wire  _T_3146; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21234.4]
  wire  _T_3148; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21236.4]
  wire  _T_3149; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21237.4]
  wire  _T_3160; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21254.4]
  wire  _T_3161; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21255.4]
  wire  _T_3163; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21257.4]
  wire  _T_3165; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21259.4]
  wire [1:0] _T_3166; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21260.4]
  wire [1:0] _T_3167; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21261.4]
  wire  _T_3168; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21262.4]
  wire  _T_3169; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21264.4]
  wire  _T_3171; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21266.4]
  wire  _T_3173; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21268.4]
  wire  _T_3174; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21269.4]
  wire  _T_3175; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21274.4]
  wire  _T_3176; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21275.4]
  wire  _T_3177; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21276.4]
  wire  _T_3179; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21278.4]
  wire  _T_3180; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21279.4]
  wire  _T_3191; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21296.4]
  wire  _T_3192; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21297.4]
  wire  _T_3194; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21299.4]
  wire  _T_3196; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21301.4]
  wire [1:0] _T_3197; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21302.4]
  wire [1:0] _T_3198; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21303.4]
  wire  _T_3199; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21304.4]
  wire  _T_3200; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21306.4]
  wire  _T_3202; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21308.4]
  wire  _T_3204; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21310.4]
  wire  _T_3205; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21311.4]
  wire  _T_3206; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21316.4]
  wire  _T_3207; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21317.4]
  wire  _T_3208; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21318.4]
  wire  _T_3210; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21320.4]
  wire  _T_3211; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21321.4]
  wire  _T_3222; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21338.4]
  wire  _T_3223; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21339.4]
  wire  _T_3225; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21341.4]
  wire  _T_3227; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21343.4]
  wire [1:0] _T_3228; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21344.4]
  wire [1:0] _T_3229; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21345.4]
  wire  _T_3230; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21346.4]
  wire  _T_3231; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21348.4]
  wire  _T_3233; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21350.4]
  wire  _T_3235; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21352.4]
  wire  _T_3236; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21353.4]
  wire  _T_3237; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21358.4]
  wire  _T_3238; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21359.4]
  wire  _T_3239; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21360.4]
  wire  _T_3241; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21362.4]
  wire  _T_3242; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21363.4]
  wire  _T_3253; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21380.4]
  wire  _T_3254; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21381.4]
  wire  _T_3256; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21383.4]
  wire  _T_3258; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21385.4]
  wire [1:0] _T_3259; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21386.4]
  wire [1:0] _T_3260; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21387.4]
  wire  _T_3261; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21388.4]
  wire  _T_3262; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21390.4]
  wire  _T_3264; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21392.4]
  wire  _T_3266; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21394.4]
  wire  _T_3267; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21395.4]
  wire  _T_3268; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21400.4]
  wire  _T_3269; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21401.4]
  wire  _T_3270; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21402.4]
  wire  _T_3272; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21404.4]
  wire  _T_3273; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21405.4]
  wire  _T_3284; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21422.4]
  wire  _T_3285; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21423.4]
  wire  _T_3287; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21425.4]
  wire  _T_3289; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21427.4]
  wire [1:0] _T_3290; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21428.4]
  wire [1:0] _T_3291; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21429.4]
  wire  _T_3292; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21430.4]
  wire  _T_3293; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21432.4]
  wire  _T_3295; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21434.4]
  wire  _T_3297; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21436.4]
  wire  _T_3298; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21437.4]
  wire  _T_3299; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21442.4]
  wire  _T_3300; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21443.4]
  wire  _T_3301; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21444.4]
  wire  _T_3303; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21446.4]
  wire  _T_3304; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21447.4]
  wire  _T_3315; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21464.4]
  wire  _T_3316; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21465.4]
  wire  _T_3318; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21467.4]
  wire  _T_3320; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21469.4]
  wire [1:0] _T_3321; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21470.4]
  wire [1:0] _T_3322; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21471.4]
  wire  _T_3323; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21472.4]
  wire  _T_3324; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21474.4]
  wire  _T_3326; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21476.4]
  wire  _T_3328; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21478.4]
  wire  _T_3329; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21479.4]
  wire  _T_3330; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21484.4]
  wire  _T_3331; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21485.4]
  wire  _T_3332; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21486.4]
  wire  _T_3334; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21488.4]
  wire  _T_3335; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21489.4]
  wire  _T_3346; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21506.4]
  wire  _T_3347; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21507.4]
  wire  _T_3349; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21509.4]
  wire  _T_3351; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21511.4]
  wire [1:0] _T_3352; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21512.4]
  wire [1:0] _T_3353; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21513.4]
  wire  _T_3354; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21514.4]
  wire  _T_3355; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21516.4]
  wire  _T_3357; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21518.4]
  wire  _T_3359; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21520.4]
  wire  _T_3360; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21521.4]
  wire  _T_3361; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21526.4]
  wire  _T_3362; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21527.4]
  wire  _T_3363; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21528.4]
  wire  _T_3365; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21530.4]
  wire  _T_3366; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21531.4]
  wire  _T_3377; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21548.4]
  wire  _T_3378; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21549.4]
  wire  _T_3380; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21551.4]
  wire  _T_3382; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21553.4]
  wire [1:0] _T_3383; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21554.4]
  wire [1:0] _T_3384; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21555.4]
  wire  _T_3385; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21556.4]
  wire  _T_3386; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21558.4]
  wire  _T_3388; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21560.4]
  wire  _T_3390; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21562.4]
  wire  _T_3391; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21563.4]
  wire  _T_3392; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21568.4]
  wire  _T_3393; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21569.4]
  wire  _T_3394; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21570.4]
  wire  _T_3396; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21572.4]
  wire  _T_3397; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21573.4]
  wire  _T_3408; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21590.4]
  wire  _T_3409; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21591.4]
  wire  _T_3411; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21593.4]
  wire  _T_3413; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21595.4]
  wire [1:0] _T_3414; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21596.4]
  wire [1:0] _T_3415; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21597.4]
  wire  _T_3416; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21598.4]
  wire  _T_3417; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21600.4]
  wire  _T_3419; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21602.4]
  wire  _T_3421; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21604.4]
  wire  _T_3422; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21605.4]
  wire  _T_3423; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21610.4]
  wire  _T_3424; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21611.4]
  wire  _T_3425; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21612.4]
  wire  _T_3427; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21614.4]
  wire  _T_3428; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21615.4]
  wire  _T_3439; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21632.4]
  wire  _T_3440; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21633.4]
  wire  _T_3442; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21635.4]
  wire  _T_3444; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21637.4]
  wire [1:0] _T_3445; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21638.4]
  wire [1:0] _T_3446; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21639.4]
  wire  _T_3447; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21640.4]
  wire  _T_3448; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21642.4]
  wire  _T_3450; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21644.4]
  wire  _T_3452; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21646.4]
  wire  _T_3453; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21647.4]
  wire  _T_3454; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21652.4]
  wire  _T_3455; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21653.4]
  wire  _T_3456; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21654.4]
  wire  _T_3458; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21656.4]
  wire  _T_3459; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21657.4]
  wire  _T_3470; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21674.4]
  wire  _T_3471; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21675.4]
  wire  _T_3473; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21677.4]
  wire  _T_3475; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21679.4]
  wire [1:0] _T_3476; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21680.4]
  wire [1:0] _T_3477; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21681.4]
  wire  _T_3478; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21682.4]
  wire  _T_3479; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21684.4]
  wire  _T_3481; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21686.4]
  wire  _T_3483; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21688.4]
  wire  _T_3484; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21689.4]
  wire  _T_3485; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21694.4]
  wire  _T_3486; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21695.4]
  wire  _T_3487; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21696.4]
  wire  _T_3489; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21698.4]
  wire  _T_3490; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21699.4]
  wire  _T_3501; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21716.4]
  wire  _T_3502; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21717.4]
  wire  _T_3504; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21719.4]
  wire  _T_3506; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21721.4]
  wire [1:0] _T_3507; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21722.4]
  wire [1:0] _T_3508; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21723.4]
  wire  _T_3509; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21724.4]
  wire  _T_3510; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21726.4]
  wire  _T_3512; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21728.4]
  wire  _T_3514; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21730.4]
  wire  _T_3515; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21731.4]
  wire  _T_3516; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21736.4]
  wire  _T_3517; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21737.4]
  wire  _T_3518; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21738.4]
  wire  _T_3520; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21740.4]
  wire  _T_3521; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21741.4]
  wire  _T_3532; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21758.4]
  wire  _T_3533; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21759.4]
  wire  _T_3535; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21761.4]
  wire  _T_3537; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21763.4]
  wire [1:0] _T_3538; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21764.4]
  wire [1:0] _T_3539; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21765.4]
  wire  _T_3540; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21766.4]
  wire  _T_3541; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21768.4]
  wire  _T_3543; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21770.4]
  wire  _T_3545; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21772.4]
  wire  _T_3546; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21773.4]
  wire  _T_3547; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21778.4]
  wire  _T_3548; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21779.4]
  wire  _T_3549; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21780.4]
  wire  _T_3551; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21782.4]
  wire  _T_3552; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21783.4]
  wire  _T_3563; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21800.4]
  wire  _T_3564; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21801.4]
  wire  _T_3566; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21803.4]
  wire  _T_3568; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21805.4]
  wire [1:0] _T_3569; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21806.4]
  wire [1:0] _T_3570; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21807.4]
  wire  _T_3571; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21808.4]
  wire  _T_3572; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21810.4]
  wire  _T_3574; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21812.4]
  wire  _T_3576; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21814.4]
  wire  _T_3577; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21815.4]
  wire  _T_3578; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21820.4]
  wire  _T_3579; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21821.4]
  wire  _T_3580; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21822.4]
  wire  _T_3582; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21824.4]
  wire  _T_3583; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21825.4]
  wire  _T_3594; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21842.4]
  wire  _T_3595; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21843.4]
  wire  _T_3597; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21845.4]
  wire  _T_3599; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21847.4]
  wire [1:0] _T_3600; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21848.4]
  wire [1:0] _T_3601; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21849.4]
  wire  _T_3602; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21850.4]
  wire  _T_3603; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21852.4]
  wire  _T_3605; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21854.4]
  wire  _T_3607; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21856.4]
  wire  _T_3608; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21857.4]
  wire  _T_3609; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21862.4]
  wire  _T_3610; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21863.4]
  wire  _T_3611; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21864.4]
  wire  _T_3613; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21866.4]
  wire  _T_3614; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21867.4]
  wire  _T_3625; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21884.4]
  wire  _T_3626; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21885.4]
  wire  _T_3628; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21887.4]
  wire  _T_3630; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21889.4]
  wire [1:0] _T_3631; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21890.4]
  wire [1:0] _T_3632; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21891.4]
  wire  _T_3633; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21892.4]
  wire  _T_3634; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21894.4]
  wire  _T_3636; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21896.4]
  wire  _T_3638; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21898.4]
  wire  _T_3639; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21899.4]
  wire  _T_3640; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21904.4]
  wire  _T_3641; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21905.4]
  wire  _T_3642; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21906.4]
  wire  _T_3644; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21908.4]
  wire  _T_3645; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21909.4]
  wire  _T_3656; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21926.4]
  wire  _T_3657; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21927.4]
  wire  _T_3659; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21929.4]
  wire  _T_3661; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21931.4]
  wire [1:0] _T_3662; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21932.4]
  wire [1:0] _T_3663; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21933.4]
  wire  _T_3664; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21934.4]
  wire  _T_3665; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21936.4]
  wire  _T_3667; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21938.4]
  wire  _T_3669; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21940.4]
  wire  _T_3670; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21941.4]
  wire  _T_3671; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21946.4]
  wire  _T_3672; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21947.4]
  wire  _T_3673; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21948.4]
  wire  _T_3675; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21950.4]
  wire  _T_3676; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21951.4]
  wire  _T_3687; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21968.4]
  wire  _T_3688; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21969.4]
  wire  _T_3690; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21971.4]
  wire  _T_3692; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21973.4]
  wire [1:0] _T_3693; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21974.4]
  wire [1:0] _T_3694; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21975.4]
  wire  _T_3695; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21976.4]
  wire  _T_3696; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21978.4]
  wire  _T_3698; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21980.4]
  wire  _T_3700; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21982.4]
  wire  _T_3701; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21983.4]
  wire  _T_3702; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21988.4]
  wire  _T_3703; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21989.4]
  wire  _T_3704; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21990.4]
  wire  _T_3706; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21992.4]
  wire  _T_3707; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21993.4]
  wire  _T_3718; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22010.4]
  wire  _T_3719; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22011.4]
  wire  _T_3721; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22013.4]
  wire  _T_3723; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22015.4]
  wire [1:0] _T_3724; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22016.4]
  wire [1:0] _T_3725; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22017.4]
  wire  _T_3726; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22018.4]
  wire  _T_3727; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22020.4]
  wire  _T_3729; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22022.4]
  wire  _T_3731; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22024.4]
  wire  _T_3732; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22025.4]
  wire  _T_3733; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22030.4]
  wire  _T_3734; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22031.4]
  wire  _T_3735; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22032.4]
  wire  _T_3737; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22034.4]
  wire  _T_3738; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22035.4]
  wire  _T_3749; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22052.4]
  wire  _T_3750; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22053.4]
  wire  _T_3752; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22055.4]
  wire  _T_3754; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22057.4]
  wire [1:0] _T_3755; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22058.4]
  wire [1:0] _T_3756; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22059.4]
  wire  _T_3757; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22060.4]
  wire  _T_3758; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22062.4]
  wire  _T_3760; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22064.4]
  wire  _T_3762; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22066.4]
  wire  _T_3763; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22067.4]
  wire  _T_3764; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22072.4]
  wire  _T_3765; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22073.4]
  wire  _T_3766; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22074.4]
  wire  _T_3768; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22076.4]
  wire  _T_3769; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22077.4]
  wire  _T_3780; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22094.4]
  wire  _T_3781; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22095.4]
  wire  _T_3783; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22097.4]
  wire  _T_3785; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22099.4]
  wire [1:0] _T_3786; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22100.4]
  wire [1:0] _T_3787; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22101.4]
  wire  _T_3788; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22102.4]
  wire  _T_3789; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22104.4]
  wire  _T_3791; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22106.4]
  wire  _T_3793; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22108.4]
  wire  _T_3794; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22109.4]
  wire  _T_3795; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22114.4]
  wire  _T_3796; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22115.4]
  wire  _T_3797; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22116.4]
  wire  _T_3799; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22118.4]
  wire  _T_3800; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22119.4]
  wire  _T_3811; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22136.4]
  wire  _T_3812; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22137.4]
  wire  _T_3814; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22139.4]
  wire  _T_3816; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22141.4]
  wire [1:0] _T_3817; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22142.4]
  wire [1:0] _T_3818; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22143.4]
  wire  _T_3819; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22144.4]
  wire  _T_3820; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22146.4]
  wire  _T_3822; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22148.4]
  wire  _T_3824; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22150.4]
  wire  _T_3825; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22151.4]
  wire  _T_3826; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22156.4]
  wire  _T_3827; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22157.4]
  wire  _T_3828; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22158.4]
  wire  _T_3830; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22160.4]
  wire  _T_3831; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22161.4]
  wire  _T_3842; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22178.4]
  wire  _T_3843; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22179.4]
  wire  _T_3845; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22181.4]
  wire  _T_3847; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22183.4]
  wire [1:0] _T_3848; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22184.4]
  wire [1:0] _T_3849; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22185.4]
  wire  _T_3850; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22186.4]
  wire  _T_3851; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22188.4]
  wire  _T_3853; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22190.4]
  wire  _T_3855; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22192.4]
  wire  _T_3856; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22193.4]
  wire  _T_3857; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22198.4]
  wire  _T_3858; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22199.4]
  wire  _T_3859; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22200.4]
  wire  _T_3861; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22202.4]
  wire  _T_3862; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22203.4]
  wire  _T_3873; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22220.4]
  wire  _T_3874; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22221.4]
  wire  _T_3876; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22223.4]
  wire  _T_3878; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22225.4]
  wire [1:0] _T_3879; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22226.4]
  wire [1:0] _T_3880; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22227.4]
  wire  _T_3881; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22228.4]
  wire  _T_3882; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22230.4]
  wire  _T_3884; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22232.4]
  wire  _T_3886; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22234.4]
  wire  _T_3887; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22235.4]
  wire  _T_3888; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22240.4]
  wire  _T_3889; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22241.4]
  wire  _T_3890; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22242.4]
  wire  _T_3892; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22244.4]
  wire  _T_3893; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22245.4]
  wire  _T_3904; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22262.4]
  wire  _T_3905; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22263.4]
  wire  _T_3907; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22265.4]
  wire  _T_3909; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22267.4]
  wire [1:0] _T_3910; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22268.4]
  wire [1:0] _T_3911; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22269.4]
  wire  _T_3912; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22270.4]
  wire  _T_3913; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22272.4]
  wire  _T_3915; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22274.4]
  wire  _T_3917; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22276.4]
  wire  _T_3918; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22277.4]
  wire  _T_3919; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22282.4]
  wire  _T_3920; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22283.4]
  wire  _T_3921; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22284.4]
  wire  _T_3923; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22286.4]
  wire  _T_3924; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22287.4]
  wire  _T_3935; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22304.4]
  wire  _T_3936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22305.4]
  wire  _T_3938; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22307.4]
  wire  _T_3940; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22309.4]
  wire [1:0] _T_3941; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22310.4]
  wire [1:0] _T_3942; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22311.4]
  wire  _T_3943; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22312.4]
  wire  _T_3944; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22314.4]
  wire  _T_3946; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22316.4]
  wire  _T_3948; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22318.4]
  wire  _T_3949; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22319.4]
  wire  _T_3950; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22324.4]
  wire  _T_3951; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22325.4]
  wire  _T_3952; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22326.4]
  wire  _T_3954; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22328.4]
  wire  _T_3955; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22329.4]
  wire  _T_3966; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22346.4]
  wire  _T_3967; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22347.4]
  wire  _T_3969; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22349.4]
  wire  _T_3971; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22351.4]
  wire [1:0] _T_3972; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22352.4]
  wire [1:0] _T_3973; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22353.4]
  wire  _T_3974; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22354.4]
  wire  _T_3975; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22356.4]
  wire  _T_3977; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22358.4]
  wire  _T_3979; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22360.4]
  wire  _T_3980; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22361.4]
  wire  _T_3981; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22366.4]
  wire  _T_3982; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22367.4]
  wire  _T_3983; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22368.4]
  wire  _T_3985; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22370.4]
  wire  _T_3986; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22371.4]
  wire  _T_3997; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22388.4]
  wire  _T_3998; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22389.4]
  wire  _T_4000; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22391.4]
  wire  _T_4002; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22393.4]
  wire [1:0] _T_4003; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22394.4]
  wire [1:0] _T_4004; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22395.4]
  wire  _T_4005; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22396.4]
  wire  _T_4006; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22398.4]
  wire  _T_4008; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22400.4]
  wire  _T_4010; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22402.4]
  wire  _T_4011; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22403.4]
  wire  _T_4012; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22408.4]
  wire  _T_4013; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22409.4]
  wire  _T_4014; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22410.4]
  wire  _T_4016; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22412.4]
  wire  _T_4017; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22413.4]
  wire  _T_4028; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22430.4]
  wire  _T_4029; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22431.4]
  wire  _T_4031; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22433.4]
  wire  _T_4033; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22435.4]
  wire [1:0] _T_4034; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22436.4]
  wire [1:0] _T_4035; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22437.4]
  wire  _T_4036; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22438.4]
  wire  _T_4037; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22440.4]
  wire  _T_4039; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22442.4]
  wire  _T_4041; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22444.4]
  wire  _T_4042; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22445.4]
  wire  _T_4043; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22450.4]
  wire  _T_4044; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22451.4]
  wire  _T_4045; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22452.4]
  wire  _T_4047; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22454.4]
  wire  _T_4048; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22455.4]
  wire  _T_4059; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22472.4]
  wire  _T_4060; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22473.4]
  wire  _T_4062; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22475.4]
  wire  _T_4064; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22477.4]
  wire [1:0] _T_4065; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22478.4]
  wire [1:0] _T_4066; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22479.4]
  wire  _T_4067; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22480.4]
  wire  _T_4068; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22482.4]
  wire  _T_4070; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22484.4]
  wire  _T_4072; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22486.4]
  wire  _T_4073; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22487.4]
  wire  _T_4074; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22492.4]
  wire  _T_4075; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22493.4]
  wire  _T_4076; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22494.4]
  wire  _T_4078; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22496.4]
  wire  _T_4079; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22497.4]
  wire  _T_4090; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22514.4]
  wire  _T_4091; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22515.4]
  wire  _T_4093; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22517.4]
  wire  _T_4095; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22519.4]
  wire [1:0] _T_4096; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22520.4]
  wire [1:0] _T_4097; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22521.4]
  wire  _T_4098; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22522.4]
  wire  _T_4099; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22524.4]
  wire  _T_4101; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22526.4]
  wire  _T_4103; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22528.4]
  wire  _T_4104; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22529.4]
  wire  _T_4105; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22534.4]
  wire  _T_4106; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22535.4]
  wire  _T_4107; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22536.4]
  wire  _T_4109; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22538.4]
  wire  _T_4110; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22539.4]
  wire  _T_4121; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22556.4]
  wire  _T_4122; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22557.4]
  wire  _T_4124; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22559.4]
  wire  _T_4126; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22561.4]
  wire [1:0] _T_4127; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22562.4]
  wire [1:0] _T_4128; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22563.4]
  wire  _T_4129; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22564.4]
  wire  _T_4130; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22566.4]
  wire  _T_4132; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22568.4]
  wire  _T_4134; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22570.4]
  wire  _T_4135; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22571.4]
  wire  _T_4136; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22576.4]
  wire  _T_4137; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22577.4]
  wire  _T_4138; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22578.4]
  wire  _T_4140; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22580.4]
  wire  _T_4141; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22581.4]
  wire  _T_4152; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22598.4]
  wire  _T_4153; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22599.4]
  wire  _T_4155; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22601.4]
  wire  _T_4157; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22603.4]
  wire [1:0] _T_4158; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22604.4]
  wire [1:0] _T_4159; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22605.4]
  wire  _T_4160; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22606.4]
  wire  _T_4161; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22608.4]
  wire  _T_4163; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22610.4]
  wire  _T_4165; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22612.4]
  wire  _T_4166; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22613.4]
  wire  _T_4167; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22618.4]
  wire  _T_4168; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22619.4]
  wire  _T_4169; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22620.4]
  wire  _T_4171; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22622.4]
  wire  _T_4172; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22623.4]
  wire  _T_4183; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22640.4]
  wire  _T_4184; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22641.4]
  wire  _T_4186; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22643.4]
  wire  _T_4188; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22645.4]
  wire [1:0] _T_4189; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22646.4]
  wire [1:0] _T_4190; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22647.4]
  wire  _T_4191; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22648.4]
  wire  _T_4192; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22650.4]
  wire  _T_4194; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22652.4]
  wire  _T_4196; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22654.4]
  wire  _T_4197; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22655.4]
  wire  _T_4198; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22660.4]
  wire  _T_4199; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22661.4]
  wire  _T_4200; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22662.4]
  wire  _T_4202; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22664.4]
  wire  _T_4203; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22665.4]
  wire  _T_4214; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22682.4]
  wire  _T_4215; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22683.4]
  wire  _T_4217; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22685.4]
  wire  _T_4219; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22687.4]
  wire [1:0] _T_4220; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22688.4]
  wire [1:0] _T_4221; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22689.4]
  wire  _T_4222; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22690.4]
  wire  _T_4223; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22692.4]
  wire  _T_4225; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22694.4]
  wire  _T_4227; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22696.4]
  wire  _T_4228; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22697.4]
  wire  _T_4229; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22702.4]
  wire  _T_4230; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22703.4]
  wire  _T_4231; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22704.4]
  wire  _T_4233; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22706.4]
  wire  _T_4234; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22707.4]
  wire  _T_4245; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22724.4]
  wire  _T_4246; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22725.4]
  wire  _T_4248; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22727.4]
  wire  _T_4250; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22729.4]
  wire [1:0] _T_4251; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22730.4]
  wire [1:0] _T_4252; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22731.4]
  wire  _T_4253; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22732.4]
  wire  _T_4254; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22734.4]
  wire  _T_4256; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22736.4]
  wire  _T_4258; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22738.4]
  wire  _T_4259; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22739.4]
  wire  _T_4260; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22744.4]
  wire  _T_4261; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22745.4]
  wire  _T_4262; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22746.4]
  wire  _T_4264; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22748.4]
  wire  _T_4265; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22749.4]
  wire  _T_4276; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22766.4]
  wire  _T_4277; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22767.4]
  wire  _T_4279; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22769.4]
  wire  _T_4281; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22771.4]
  wire [1:0] _T_4282; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22772.4]
  wire [1:0] _T_4283; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22773.4]
  wire  _T_4284; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22774.4]
  wire  _T_4285; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22776.4]
  wire  _T_4287; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22778.4]
  wire  _T_4289; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22780.4]
  wire  _T_4290; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22781.4]
  wire  _T_4291; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22786.4]
  wire  _T_4292; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22787.4]
  wire  _T_4293; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22788.4]
  wire  _T_4295; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22790.4]
  wire  _T_4296; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22791.4]
  wire  _T_4307; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22808.4]
  wire  _T_4308; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22809.4]
  wire  _T_4310; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22811.4]
  wire  _T_4312; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22813.4]
  wire [1:0] _T_4313; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22814.4]
  wire [1:0] _T_4314; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22815.4]
  wire  _T_4315; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22816.4]
  wire  _T_4316; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22818.4]
  wire  _T_4318; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22820.4]
  wire  _T_4320; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22822.4]
  wire  _T_4321; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22823.4]
  wire  _T_4322; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22828.4]
  wire  _T_4323; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22829.4]
  wire  _T_4324; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22830.4]
  wire  _T_4326; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22832.4]
  wire  _T_4327; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22833.4]
  wire  _T_4338; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22850.4]
  wire  _T_4339; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22851.4]
  wire  _T_4341; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22853.4]
  wire  _T_4343; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22855.4]
  wire [1:0] _T_4344; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22856.4]
  wire [1:0] _T_4345; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22857.4]
  wire  _T_4346; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22858.4]
  wire  _T_4347; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22860.4]
  wire  _T_4349; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22862.4]
  wire  _T_4351; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22864.4]
  wire  _T_4352; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22865.4]
  wire  _T_4353; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22870.4]
  wire  _T_4354; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22871.4]
  wire  _T_4355; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22872.4]
  wire  _T_4357; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22874.4]
  wire  _T_4358; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22875.4]
  wire  _T_4369; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22892.4]
  wire  _T_4370; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22893.4]
  wire  _T_4372; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22895.4]
  wire  _T_4374; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22897.4]
  wire [1:0] _T_4375; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22898.4]
  wire [1:0] _T_4376; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22899.4]
  wire  _T_4377; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22900.4]
  wire  _T_4378; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22902.4]
  wire  _T_4380; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22904.4]
  wire  _T_4382; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22906.4]
  wire  _T_4383; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22907.4]
  wire  _T_4384; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22912.4]
  wire  _T_4385; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22913.4]
  wire  _T_4386; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22914.4]
  wire  _T_4388; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22916.4]
  wire  _T_4389; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22917.4]
  wire  _T_4400; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22934.4]
  wire  _T_4401; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22935.4]
  wire  _T_4403; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22937.4]
  wire  _T_4405; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22939.4]
  wire [1:0] _T_4406; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22940.4]
  wire [1:0] _T_4407; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22941.4]
  wire  _T_4408; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22942.4]
  wire  _T_4409; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22944.4]
  wire  _T_4411; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22946.4]
  wire  _T_4413; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22948.4]
  wire  _T_4414; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22949.4]
  wire  _T_4415; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22954.4]
  wire  _T_4416; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22955.4]
  wire  _T_4417; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22956.4]
  wire  _T_4419; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22958.4]
  wire  _T_4420; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22959.4]
  wire  _T_4431; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22976.4]
  wire  _T_4432; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22977.4]
  wire  _T_4434; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22979.4]
  wire  _T_4436; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22981.4]
  wire [1:0] _T_4437; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22982.4]
  wire [1:0] _T_4438; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22983.4]
  wire  _T_4439; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22984.4]
  wire  _T_4440; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22986.4]
  wire  _T_4442; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22988.4]
  wire  _T_4444; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22990.4]
  wire  _T_4445; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22991.4]
  wire  _T_4446; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22996.4]
  wire  _T_4447; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22997.4]
  wire  _T_4448; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22998.4]
  wire  _T_4450; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23000.4]
  wire  _T_4451; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23001.4]
  wire  _T_4462; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23018.4]
  wire  _T_4463; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23019.4]
  wire  _T_4465; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23021.4]
  wire  _T_4467; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23023.4]
  wire [1:0] _T_4468; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23024.4]
  wire [1:0] _T_4469; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23025.4]
  wire  _T_4470; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23026.4]
  wire  _T_4471; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23028.4]
  wire  _T_4473; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23030.4]
  wire  _T_4475; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23032.4]
  wire  _T_4476; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23033.4]
  wire  _T_4477; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23038.4]
  wire  _T_4478; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23039.4]
  wire  _T_4479; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23040.4]
  wire  _T_4481; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23042.4]
  wire  _T_4482; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23043.4]
  wire  _T_4493; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23060.4]
  wire  _T_4494; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23061.4]
  wire  _T_4496; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23063.4]
  wire  _T_4498; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23065.4]
  wire [1:0] _T_4499; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23066.4]
  wire [1:0] _T_4500; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23067.4]
  wire  _T_4501; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23068.4]
  wire  _T_4502; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23070.4]
  wire  _T_4504; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23072.4]
  wire  _T_4506; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23074.4]
  wire  _T_4507; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23075.4]
  wire  _T_4508; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23080.4]
  wire  _T_4509; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23081.4]
  wire  _T_4510; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23082.4]
  wire  _T_4512; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23084.4]
  wire  _T_4513; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23085.4]
  wire  _T_4524; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23102.4]
  wire  _T_4525; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23103.4]
  wire  _T_4527; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23105.4]
  wire  _T_4529; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23107.4]
  wire [1:0] _T_4530; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23108.4]
  wire [1:0] _T_4531; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23109.4]
  wire  _T_4532; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23110.4]
  wire  _T_4533; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23112.4]
  wire  _T_4535; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23114.4]
  wire  _T_4537; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23116.4]
  wire  _T_4538; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23117.4]
  wire  _T_4539; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23122.4]
  wire  _T_4540; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23123.4]
  wire  _T_4541; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23124.4]
  wire  _T_4543; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23126.4]
  wire  _T_4544; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23127.4]
  wire  _T_4555; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23144.4]
  wire  _T_4556; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23145.4]
  wire  _T_4558; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23147.4]
  wire  _T_4560; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23149.4]
  wire [1:0] _T_4561; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23150.4]
  wire [1:0] _T_4562; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23151.4]
  wire  _T_4563; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23152.4]
  wire  _T_4564; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23154.4]
  wire  _T_4566; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23156.4]
  wire  _T_4568; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23158.4]
  wire  _T_4569; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23159.4]
  wire  _T_4570; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23164.4]
  wire  _T_4571; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23165.4]
  wire  _T_4572; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23166.4]
  wire  _T_4574; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23168.4]
  wire  _T_4575; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23169.4]
  wire  _T_4586; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23186.4]
  wire  _T_4587; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23187.4]
  wire  _T_4589; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23189.4]
  wire  _T_4591; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23191.4]
  wire [1:0] _T_4592; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23192.4]
  wire [1:0] _T_4593; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23193.4]
  wire  _T_4594; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23194.4]
  wire  _T_4595; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23196.4]
  wire  _T_4597; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23198.4]
  wire  _T_4599; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23200.4]
  wire  _T_4600; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23201.4]
  wire  _T_4601; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23206.4]
  wire  _T_4602; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23207.4]
  wire  _T_4603; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23208.4]
  wire  _T_4605; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23210.4]
  wire  _T_4606; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23211.4]
  wire  _T_4617; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23228.4]
  wire  _T_4618; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23229.4]
  wire  _T_4620; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23231.4]
  wire  _T_4622; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23233.4]
  wire [1:0] _T_4623; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23234.4]
  wire [1:0] _T_4624; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23235.4]
  wire  _T_4625; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23236.4]
  wire  _T_4626; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23238.4]
  wire  _T_4628; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23240.4]
  wire  _T_4630; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23242.4]
  wire  _T_4631; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23243.4]
  wire  _T_4632; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23248.4]
  wire  _T_4633; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23249.4]
  wire  _T_4634; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23250.4]
  wire  _T_4636; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23252.4]
  wire  _T_4637; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23253.4]
  wire  _T_4648; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23270.4]
  wire  _T_4649; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23271.4]
  wire  _T_4651; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23273.4]
  wire  _T_4653; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23275.4]
  wire [1:0] _T_4654; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23276.4]
  wire [1:0] _T_4655; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23277.4]
  wire  _T_4656; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23278.4]
  wire  _T_4657; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23280.4]
  wire  _T_4659; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23282.4]
  wire  _T_4661; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23284.4]
  wire  _T_4662; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23285.4]
  wire  _T_4663; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23290.4]
  wire  _T_4664; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23291.4]
  wire  _T_4665; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23292.4]
  wire  _T_4667; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23294.4]
  wire  _T_4668; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23295.4]
  wire  _T_4679; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23312.4]
  wire  _T_4680; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23313.4]
  wire  _T_4682; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23315.4]
  wire  _T_4684; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23317.4]
  wire [1:0] _T_4685; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23318.4]
  wire [1:0] _T_4686; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23319.4]
  wire  _T_4687; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23320.4]
  wire  _T_4688; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23322.4]
  wire  _T_4690; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23324.4]
  wire  _T_4692; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23326.4]
  wire  _T_4693; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23327.4]
  wire  _T_4694; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23332.4]
  wire  _T_4695; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23333.4]
  wire  _T_4696; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23334.4]
  wire  _T_4698; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23336.4]
  wire  _T_4699; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23337.4]
  wire  _T_4710; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23354.4]
  wire  _T_4711; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23355.4]
  wire  _T_4713; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23357.4]
  wire  _T_4715; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23359.4]
  wire [1:0] _T_4716; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23360.4]
  wire [1:0] _T_4717; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23361.4]
  wire  _T_4718; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23362.4]
  wire  _T_4719; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23364.4]
  wire  _T_4721; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23366.4]
  wire  _T_4723; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23368.4]
  wire  _T_4724; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23369.4]
  wire  _T_4725; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23374.4]
  wire  _T_4726; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23375.4]
  wire  _T_4727; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23376.4]
  wire  _T_4729; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23378.4]
  wire  _T_4730; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23379.4]
  wire  _T_4741; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23396.4]
  wire  _T_4742; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23397.4]
  wire  _T_4744; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23399.4]
  wire  _T_4746; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23401.4]
  wire [1:0] _T_4747; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23402.4]
  wire [1:0] _T_4748; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23403.4]
  wire  _T_4749; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23404.4]
  wire  _T_4750; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23406.4]
  wire  _T_4752; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23408.4]
  wire  _T_4754; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23410.4]
  wire  _T_4755; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23411.4]
  wire  _T_4756; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23416.4]
  wire  _T_4757; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23417.4]
  wire  _T_4758; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23418.4]
  wire  _T_4760; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23420.4]
  wire  _T_4761; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23421.4]
  wire  _T_4772; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23438.4]
  wire  _T_4773; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23439.4]
  wire  _T_4775; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23441.4]
  wire  _T_4777; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23443.4]
  wire [1:0] _T_4778; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23444.4]
  wire [1:0] _T_4779; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23445.4]
  wire  _T_4780; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23446.4]
  wire  _T_4781; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23448.4]
  wire  _T_4783; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23450.4]
  wire  _T_4785; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23452.4]
  wire  _T_4786; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23453.4]
  wire  _T_4787; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23458.4]
  wire  _T_4788; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23459.4]
  wire  _T_4789; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23460.4]
  wire  _T_4791; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23462.4]
  wire  _T_4792; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23463.4]
  wire  _T_4803; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23480.4]
  wire  _T_4804; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23481.4]
  wire  _T_4806; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23483.4]
  wire  _T_4808; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23485.4]
  wire [1:0] _T_4809; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23486.4]
  wire [1:0] _T_4810; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23487.4]
  wire  _T_4811; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23488.4]
  wire  _T_4812; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23490.4]
  wire  _T_4814; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23492.4]
  wire  _T_4816; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23494.4]
  wire  _T_4817; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23495.4]
  wire  _T_4818; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23500.4]
  wire  _T_4819; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23501.4]
  wire  _T_4820; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23502.4]
  wire  _T_4822; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23504.4]
  wire  _T_4823; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23505.4]
  wire  _T_4834; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23522.4]
  wire  _T_4835; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23523.4]
  wire  _T_4837; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23525.4]
  wire  _T_4839; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23527.4]
  wire [1:0] _T_4840; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23528.4]
  wire [1:0] _T_4841; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23529.4]
  wire  _T_4842; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23530.4]
  wire  _T_4843; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23532.4]
  wire  _T_4845; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23534.4]
  wire  _T_4847; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23536.4]
  wire  _T_4848; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23537.4]
  wire  _T_4849; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23542.4]
  wire  _T_4850; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23543.4]
  wire  _T_4851; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23544.4]
  wire  _T_4853; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23546.4]
  wire  _T_4854; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23547.4]
  wire  _T_4865; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23564.4]
  wire  _T_4866; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23565.4]
  wire  _T_4868; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23567.4]
  wire  _T_4870; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23569.4]
  wire [1:0] _T_4871; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23570.4]
  wire [1:0] _T_4872; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23571.4]
  wire  _T_4873; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23572.4]
  wire  _T_4874; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23574.4]
  wire  _T_4876; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23576.4]
  wire  _T_4878; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23578.4]
  wire  _T_4879; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23579.4]
  wire  _T_4880; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23584.4]
  wire  _T_4881; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23585.4]
  wire  _T_4882; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23586.4]
  wire  _T_4884; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23588.4]
  wire  _T_4885; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23589.4]
  wire  _T_4896; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23606.4]
  wire  _T_4897; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23607.4]
  wire  _T_4899; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23609.4]
  wire  _T_4901; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23611.4]
  wire [1:0] _T_4902; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23612.4]
  wire [1:0] _T_4903; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23613.4]
  wire  _T_4904; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23614.4]
  wire  _T_4905; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23616.4]
  wire  _T_4907; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23618.4]
  wire  _T_4909; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23620.4]
  wire  _T_4910; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23621.4]
  wire  _T_4911; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23626.4]
  wire  _T_4912; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23627.4]
  wire  _T_4913; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23628.4]
  wire  _T_4915; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23630.4]
  wire  _T_4916; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23631.4]
  wire  _T_4927; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23648.4]
  wire  _T_4928; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23649.4]
  wire  _T_4930; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23651.4]
  wire  _T_4932; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23653.4]
  wire [1:0] _T_4933; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23654.4]
  wire [1:0] _T_4934; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23655.4]
  wire  _T_4935; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23656.4]
  wire  _T_4936; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23658.4]
  wire  _T_4938; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23660.4]
  wire  _T_4940; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23662.4]
  wire  _T_4941; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23663.4]
  wire  _T_4942; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23668.4]
  wire  _T_4943; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23669.4]
  wire  _T_4944; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23670.4]
  wire  _T_4946; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23672.4]
  wire  _T_4947; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23673.4]
  wire  _T_4958; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23690.4]
  wire  _T_4959; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23691.4]
  wire  _T_4961; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23693.4]
  wire  _T_4963; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23695.4]
  wire [1:0] _T_4964; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23696.4]
  wire [1:0] _T_4965; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23697.4]
  wire  _T_4966; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23698.4]
  wire  _T_4967; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23700.4]
  wire  _T_4969; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23702.4]
  wire  _T_4971; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23704.4]
  wire  _T_4972; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23705.4]
  wire  _T_4973; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23710.4]
  wire  _T_4974; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23711.4]
  wire  _T_4975; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23712.4]
  wire  _T_4977; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23714.4]
  wire  _T_4978; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23715.4]
  wire  _T_4989; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23732.4]
  wire  _T_4990; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23733.4]
  wire  _T_4992; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23735.4]
  wire  _T_4994; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23737.4]
  wire [1:0] _T_4995; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23738.4]
  wire [1:0] _T_4996; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23739.4]
  wire  _T_4997; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23740.4]
  wire  _T_4998; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23742.4]
  wire  _T_5000; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23744.4]
  wire  _T_5002; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23746.4]
  wire  _T_5003; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23747.4]
  wire  _T_5004; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23752.4]
  wire  _T_5005; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23753.4]
  wire  _T_5006; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23754.4]
  wire  _T_5008; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23756.4]
  wire  _T_5009; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23757.4]
  wire  _T_5020; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23774.4]
  wire  _T_5021; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23775.4]
  wire  _T_5023; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23777.4]
  wire  _T_5025; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23779.4]
  wire [1:0] _T_5026; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23780.4]
  wire [1:0] _T_5027; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23781.4]
  wire  _T_5028; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23782.4]
  wire  _T_5029; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23784.4]
  wire  _T_5031; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23786.4]
  wire  _T_5033; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23788.4]
  wire  _T_5034; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23789.4]
  wire  _T_5035; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23794.4]
  wire  _T_5036; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23795.4]
  wire  _T_5037; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23796.4]
  wire  _T_5039; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23798.4]
  wire  _T_5040; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23799.4]
  wire  _T_5051; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23816.4]
  wire  _T_5052; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23817.4]
  wire  _T_5054; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23819.4]
  wire  _T_5056; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23821.4]
  wire [1:0] _T_5057; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23822.4]
  wire [1:0] _T_5058; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23823.4]
  wire  _T_5059; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23824.4]
  wire  _T_5060; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23826.4]
  wire  _T_5062; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23828.4]
  wire  _T_5064; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23830.4]
  wire  _T_5065; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23831.4]
  wire  _T_5066; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23836.4]
  wire  _T_5067; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23837.4]
  wire  _T_5068; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23838.4]
  wire  _T_5070; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23840.4]
  wire  _T_5071; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23841.4]
  wire  _T_5082; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23858.4]
  wire  _T_5083; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23859.4]
  wire  _T_5085; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23861.4]
  wire  _T_5087; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23863.4]
  wire [1:0] _T_5088; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23864.4]
  wire [1:0] _T_5089; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23865.4]
  wire  _T_5090; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23866.4]
  wire  _T_5091; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23868.4]
  wire  _T_5093; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23870.4]
  wire  _T_5095; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23872.4]
  wire  _T_5096; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23873.4]
  wire  _T_5097; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23878.4]
  wire  _T_5098; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23879.4]
  wire  _T_5099; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23880.4]
  wire  _T_5101; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23882.4]
  wire  _T_5102; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23883.4]
  wire  _T_5113; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23900.4]
  wire  _T_5114; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23901.4]
  wire  _T_5116; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23903.4]
  wire  _T_5118; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23905.4]
  wire [1:0] _T_5119; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23906.4]
  wire [1:0] _T_5120; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23907.4]
  wire  _T_5121; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23908.4]
  wire  _T_5122; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23910.4]
  wire  _T_5124; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23912.4]
  wire  _T_5126; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23914.4]
  wire  _T_5127; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23915.4]
  wire  _T_5128; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23920.4]
  wire  _T_5129; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23921.4]
  wire  _T_5130; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23922.4]
  wire  _T_5132; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23924.4]
  wire  _T_5133; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23925.4]
  wire  _T_5144; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23942.4]
  wire  _T_5145; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23943.4]
  wire  _T_5147; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23945.4]
  wire  _T_5149; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23947.4]
  wire [1:0] _T_5150; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23948.4]
  wire [1:0] _T_5151; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23949.4]
  wire  _T_5152; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23950.4]
  wire  _T_5153; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23952.4]
  wire  _T_5155; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23954.4]
  wire  _T_5157; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23956.4]
  wire  _T_5158; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23957.4]
  wire  _T_5159; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23962.4]
  wire  _T_5160; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23963.4]
  wire  _T_5161; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23964.4]
  wire  _T_5163; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23966.4]
  wire  _T_5164; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23967.4]
  wire  _T_5175; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23984.4]
  wire  _T_5176; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23985.4]
  wire  _T_5178; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23987.4]
  wire  _T_5180; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23989.4]
  wire [1:0] _T_5181; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23990.4]
  wire [1:0] _T_5182; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23991.4]
  wire  _T_5183; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23992.4]
  wire  _T_5184; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23994.4]
  wire  _T_5186; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23996.4]
  wire  _T_5188; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23998.4]
  wire  _T_5189; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23999.4]
  wire  _T_5190; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24004.4]
  wire  _T_5191; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24005.4]
  wire  _T_5192; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24006.4]
  wire  _T_5194; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24008.4]
  wire  _T_5195; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24009.4]
  wire  _T_5206; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24026.4]
  wire  _T_5207; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24027.4]
  wire  _T_5209; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24029.4]
  wire  _T_5211; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24031.4]
  wire [1:0] _T_5212; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24032.4]
  wire [1:0] _T_5213; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24033.4]
  wire  _T_5214; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24034.4]
  wire  _T_5215; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24036.4]
  wire  _T_5217; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24038.4]
  wire  _T_5219; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24040.4]
  wire  _T_5220; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24041.4]
  wire  _T_5221; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24046.4]
  wire  _T_5222; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24047.4]
  wire  _T_5223; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24048.4]
  wire  _T_5225; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24050.4]
  wire  _T_5226; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24051.4]
  wire  _T_5237; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24068.4]
  wire  _T_5238; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24069.4]
  wire  _T_5240; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24071.4]
  wire  _T_5242; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24073.4]
  wire [1:0] _T_5243; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24074.4]
  wire [1:0] _T_5244; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24075.4]
  wire  _T_5245; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24076.4]
  wire  _T_5246; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24078.4]
  wire  _T_5248; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24080.4]
  wire  _T_5250; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24082.4]
  wire  _T_5251; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24083.4]
  wire  _T_5252; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24088.4]
  wire  _T_5253; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24089.4]
  wire  _T_5254; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24090.4]
  wire  _T_5256; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24092.4]
  wire  _T_5257; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24093.4]
  wire  _T_5268; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24110.4]
  wire  _T_5269; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24111.4]
  wire  _T_5271; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24113.4]
  wire  _T_5273; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24115.4]
  wire [1:0] _T_5274; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24116.4]
  wire [1:0] _T_5275; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24117.4]
  wire  _T_5276; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24118.4]
  wire  _T_5277; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24120.4]
  wire  _T_5279; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24122.4]
  wire  _T_5281; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24124.4]
  wire  _T_5282; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24125.4]
  wire  _T_5283; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24130.4]
  wire  _T_5284; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24131.4]
  wire  _T_5285; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24132.4]
  wire  _T_5287; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24134.4]
  wire  _T_5288; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24135.4]
  wire  _T_5299; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24152.4]
  wire  _T_5300; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24153.4]
  wire  _T_5302; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24155.4]
  wire  _T_5304; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24157.4]
  wire [1:0] _T_5305; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24158.4]
  wire [1:0] _T_5306; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24159.4]
  wire  _T_5307; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24160.4]
  wire  _T_5308; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24162.4]
  wire  _T_5310; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24164.4]
  wire  _T_5312; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24166.4]
  wire  _T_5313; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24167.4]
  wire  _T_5314; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24172.4]
  wire  _T_5315; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24173.4]
  wire  _T_5316; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24174.4]
  wire  _T_5318; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24176.4]
  wire  _T_5319; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24177.4]
  wire  _T_5330; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24194.4]
  wire  _T_5331; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24195.4]
  wire  _T_5333; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24197.4]
  wire  _T_5335; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24199.4]
  wire [1:0] _T_5336; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24200.4]
  wire [1:0] _T_5337; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24201.4]
  wire  _T_5338; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24202.4]
  wire  _T_5339; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24204.4]
  wire  _T_5341; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24206.4]
  wire  _T_5343; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24208.4]
  wire  _T_5344; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24209.4]
  wire  _T_5345; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24214.4]
  wire  _T_5346; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24215.4]
  wire  _T_5347; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24216.4]
  wire  _T_5349; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24218.4]
  wire  _T_5350; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24219.4]
  wire  _T_5361; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24236.4]
  wire  _T_5362; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24237.4]
  wire  _T_5364; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24239.4]
  wire  _T_5366; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24241.4]
  wire [1:0] _T_5367; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24242.4]
  wire [1:0] _T_5368; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24243.4]
  wire  _T_5369; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24244.4]
  wire  _T_5370; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24246.4]
  wire  _T_5372; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24248.4]
  wire  _T_5374; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24250.4]
  wire  _T_5375; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24251.4]
  wire  _T_5376; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24256.4]
  wire  _T_5377; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24257.4]
  wire  _T_5378; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24258.4]
  wire  _T_5380; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24260.4]
  wire  _T_5381; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24261.4]
  wire  _T_5392; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24278.4]
  wire  _T_5393; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24279.4]
  wire  _T_5395; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24281.4]
  wire  _T_5397; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24283.4]
  wire [1:0] _T_5398; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24284.4]
  wire [1:0] _T_5399; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24285.4]
  wire  _T_5400; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24286.4]
  wire  _T_5401; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24288.4]
  wire  _T_5403; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24290.4]
  wire  _T_5405; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24292.4]
  wire  _T_5406; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24293.4]
  wire  _T_5407; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24298.4]
  wire  _T_5408; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24299.4]
  wire  _T_5409; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24300.4]
  wire  _T_5411; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24302.4]
  wire  _T_5412; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24303.4]
  wire  _T_5423; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24320.4]
  wire  _T_5424; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24321.4]
  wire  _T_5426; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24323.4]
  wire  _T_5428; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24325.4]
  wire [1:0] _T_5429; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24326.4]
  wire [1:0] _T_5430; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24327.4]
  wire  _T_5431; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24328.4]
  wire  _T_5432; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24330.4]
  wire  _T_5434; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24332.4]
  wire  _T_5436; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24334.4]
  wire  _T_5437; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24335.4]
  wire  _T_5438; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24340.4]
  wire  _T_5439; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24341.4]
  wire  _T_5440; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24342.4]
  wire  _T_5442; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24344.4]
  wire  _T_5443; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24345.4]
  wire  _T_5454; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24362.4]
  wire  _T_5455; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24363.4]
  wire  _T_5457; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24365.4]
  wire  _T_5459; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24367.4]
  wire [1:0] _T_5460; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24368.4]
  wire [1:0] _T_5461; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24369.4]
  wire  _T_5462; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24370.4]
  wire  _T_5463; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24372.4]
  wire  _T_5465; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24374.4]
  wire  _T_5467; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24376.4]
  wire  _T_5468; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24377.4]
  wire  _T_5469; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24382.4]
  wire  _T_5470; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24383.4]
  wire  _T_5471; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24384.4]
  wire  _T_5473; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24386.4]
  wire  _T_5474; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24387.4]
  wire  _T_5485; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24404.4]
  wire  _T_5486; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24405.4]
  wire  _T_5488; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24407.4]
  wire  _T_5490; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24409.4]
  wire [1:0] _T_5491; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24410.4]
  wire [1:0] _T_5492; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24411.4]
  wire  _T_5493; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24412.4]
  wire  _T_5494; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24414.4]
  wire  _T_5496; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24416.4]
  wire  _T_5498; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24418.4]
  wire  _T_5499; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24419.4]
  wire  _T_5500; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24424.4]
  wire  _T_5501; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24425.4]
  wire  _T_5502; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24426.4]
  wire  _T_5504; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24428.4]
  wire  _T_5505; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24429.4]
  wire  _T_5516; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24446.4]
  wire  _T_5517; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24447.4]
  wire  _T_5519; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24449.4]
  wire  _T_5521; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24451.4]
  wire [1:0] _T_5522; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24452.4]
  wire [1:0] _T_5523; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24453.4]
  wire  _T_5524; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24454.4]
  wire  _T_5525; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24456.4]
  wire  _T_5527; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24458.4]
  wire  _T_5529; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24460.4]
  wire  _T_5530; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24461.4]
  wire  _T_5531; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24466.4]
  wire  _T_5532; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24467.4]
  wire  _T_5533; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24468.4]
  wire  _T_5535; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24470.4]
  wire  _T_5536; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24471.4]
  wire  _T_5547; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24488.4]
  wire  _T_5548; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24489.4]
  wire  _T_5550; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24491.4]
  wire  _T_5552; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24493.4]
  wire [1:0] _T_5553; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24494.4]
  wire [1:0] _T_5554; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24495.4]
  wire  _T_5555; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24496.4]
  wire  _T_5556; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24498.4]
  wire  _T_5558; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24500.4]
  wire  _T_5560; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24502.4]
  wire  _T_5561; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24503.4]
  wire  _T_5562; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24508.4]
  wire  _T_5563; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24509.4]
  wire  _T_5564; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24510.4]
  wire  _T_5566; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24512.4]
  wire  _T_5567; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24513.4]
  wire  _T_5578; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24530.4]
  wire  _T_5579; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24531.4]
  wire  _T_5581; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24533.4]
  wire  _T_5583; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24535.4]
  wire [1:0] _T_5584; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24536.4]
  wire [1:0] _T_5585; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24537.4]
  wire  _T_5586; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24538.4]
  wire  _T_5587; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24540.4]
  wire  _T_5589; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24542.4]
  wire  _T_5591; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24544.4]
  wire  _T_5592; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24545.4]
  wire  _T_5593; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24550.4]
  wire  _T_5594; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24551.4]
  wire  _T_5595; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24552.4]
  wire  _T_5597; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24554.4]
  wire  _T_5598; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24555.4]
  wire  _T_5609; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24572.4]
  wire  _T_5610; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24573.4]
  wire  _T_5612; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24575.4]
  wire  _T_5614; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24577.4]
  wire [1:0] _T_5615; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24578.4]
  wire [1:0] _T_5616; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24579.4]
  wire  _T_5617; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24580.4]
  wire  _T_5618; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24582.4]
  wire  _T_5620; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24584.4]
  wire  _T_5622; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24586.4]
  wire  _T_5623; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24587.4]
  wire  _T_5624; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24592.4]
  wire  _T_5625; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24593.4]
  wire  _T_5626; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24594.4]
  wire  _T_5628; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24596.4]
  wire  _T_5629; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24597.4]
  wire  _T_5640; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24614.4]
  wire  _T_5641; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24615.4]
  wire  _T_5643; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24617.4]
  wire  _T_5645; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24619.4]
  wire [1:0] _T_5646; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24620.4]
  wire [1:0] _T_5647; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24621.4]
  wire  _T_5648; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24622.4]
  wire  _T_5649; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24624.4]
  wire  _T_5651; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24626.4]
  wire  _T_5653; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24628.4]
  wire  _T_5654; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24629.4]
  wire  _T_5655; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24634.4]
  wire  _T_5656; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24635.4]
  wire  _T_5657; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24636.4]
  wire  _T_5659; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24638.4]
  wire  _T_5660; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24639.4]
  wire  _T_5671; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24656.4]
  wire  _T_5672; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24657.4]
  wire  _T_5674; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24659.4]
  wire  _T_5676; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24661.4]
  wire [1:0] _T_5677; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24662.4]
  wire [1:0] _T_5678; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24663.4]
  wire  _T_5679; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24664.4]
  wire  _T_5680; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24666.4]
  wire  _T_5682; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24668.4]
  wire  _T_5684; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24670.4]
  wire  _T_5685; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24671.4]
  wire  _T_5686; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24676.4]
  wire  _T_5687; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24677.4]
  wire  _T_5688; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24678.4]
  wire  _T_5690; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24680.4]
  wire  _T_5691; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24681.4]
  wire  _T_5702; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24698.4]
  wire  _T_5703; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24699.4]
  wire  _T_5705; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24701.4]
  wire  _T_5707; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24703.4]
  wire [1:0] _T_5708; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24704.4]
  wire [1:0] _T_5709; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24705.4]
  wire  _T_5710; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24706.4]
  wire  _T_5711; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24708.4]
  wire  _T_5713; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24710.4]
  wire  _T_5715; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24712.4]
  wire  _T_5716; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24713.4]
  wire  _T_5717; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24718.4]
  wire  _T_5718; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24719.4]
  wire  _T_5719; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24720.4]
  wire  _T_5721; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24722.4]
  wire  _T_5722; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24723.4]
  wire  _T_5733; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24740.4]
  wire  _T_5734; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24741.4]
  wire  _T_5736; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24743.4]
  wire  _T_5738; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24745.4]
  wire [1:0] _T_5739; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24746.4]
  wire [1:0] _T_5740; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24747.4]
  wire  _T_5741; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24748.4]
  wire  _T_5742; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24750.4]
  wire  _T_5744; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24752.4]
  wire  _T_5746; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24754.4]
  wire  _T_5747; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24755.4]
  wire  _T_5748; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24760.4]
  wire  _T_5749; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24761.4]
  wire  _T_5750; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24762.4]
  wire  _T_5752; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24764.4]
  wire  _T_5753; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24765.4]
  wire  _T_5764; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24782.4]
  wire  _T_5765; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24783.4]
  wire  _T_5767; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24785.4]
  wire  _T_5769; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24787.4]
  wire [1:0] _T_5770; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24788.4]
  wire [1:0] _T_5771; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24789.4]
  wire  _T_5772; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24790.4]
  wire  _T_5773; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24792.4]
  wire  _T_5775; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24794.4]
  wire  _T_5777; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24796.4]
  wire  _T_5778; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24797.4]
  wire  _T_5779; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24802.4]
  wire  _T_5780; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24803.4]
  wire  _T_5781; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24804.4]
  wire  _T_5783; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24806.4]
  wire  _T_5784; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24807.4]
  wire  _T_5795; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24824.4]
  wire  _T_5796; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24825.4]
  wire  _T_5798; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24827.4]
  wire  _T_5800; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24829.4]
  wire [1:0] _T_5801; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24830.4]
  wire [1:0] _T_5802; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24831.4]
  wire  _T_5803; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24832.4]
  wire  _T_5804; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24834.4]
  wire  _T_5806; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24836.4]
  wire  _T_5808; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24838.4]
  wire  _T_5809; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24839.4]
  wire  _T_5810; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24844.4]
  wire  _T_5811; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24845.4]
  wire  _T_5812; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24846.4]
  wire  _T_5814; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24848.4]
  wire  _T_5815; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24849.4]
  wire  _T_5826; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24866.4]
  wire  _T_5827; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24867.4]
  wire  _T_5829; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24869.4]
  wire  _T_5831; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24871.4]
  wire [1:0] _T_5832; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24872.4]
  wire [1:0] _T_5833; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24873.4]
  wire  _T_5834; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24874.4]
  wire  _T_5835; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24876.4]
  wire  _T_5837; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24878.4]
  wire  _T_5839; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24880.4]
  wire  _T_5840; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24881.4]
  wire  _T_5841; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24886.4]
  wire  _T_5842; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24887.4]
  wire  _T_5843; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24888.4]
  wire  _T_5845; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24890.4]
  wire  _T_5846; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24891.4]
  wire  _T_5857; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24908.4]
  wire  _T_5858; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24909.4]
  wire  _T_5860; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24911.4]
  wire  _T_5862; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24913.4]
  wire [1:0] _T_5863; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24914.4]
  wire [1:0] _T_5864; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24915.4]
  wire  _T_5865; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24916.4]
  wire  _T_5866; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24918.4]
  wire  _T_5868; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24920.4]
  wire  _T_5870; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24922.4]
  wire  _T_5871; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24923.4]
  wire  _T_5872; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24928.4]
  wire  _T_5873; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24929.4]
  wire  _T_5874; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24930.4]
  wire  _T_5876; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24932.4]
  wire  _T_5877; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24933.4]
  wire  _T_5888; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24950.4]
  wire  _T_5889; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24951.4]
  wire  _T_5891; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24953.4]
  wire  _T_5893; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24955.4]
  wire [1:0] _T_5894; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24956.4]
  wire [1:0] _T_5895; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24957.4]
  wire  _T_5896; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24958.4]
  wire  _T_5897; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24960.4]
  wire  _T_5899; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24962.4]
  wire  _T_5901; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24964.4]
  wire  _T_5902; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24965.4]
  wire  _T_5903; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24970.4]
  wire  _T_5904; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24971.4]
  wire  _T_5905; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24972.4]
  wire  _T_5907; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24974.4]
  wire  _T_5908; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24975.4]
  wire  _T_5919; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24992.4]
  wire  _T_5920; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24993.4]
  wire  _T_5922; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24995.4]
  wire  _T_5924; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24997.4]
  wire [1:0] _T_5925; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24998.4]
  wire [1:0] _T_5926; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24999.4]
  wire  _T_5927; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25000.4]
  wire  _T_5928; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25002.4]
  wire  _T_5930; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25004.4]
  wire  _T_5932; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25006.4]
  wire  _T_5933; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25007.4]
  wire  _T_5934; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25012.4]
  wire  _T_5935; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25013.4]
  wire  _T_5936; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25014.4]
  wire  _T_5938; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25016.4]
  wire  _T_5939; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25017.4]
  wire  _T_5950; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25034.4]
  wire  _T_5951; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25035.4]
  wire  _T_5953; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25037.4]
  wire  _T_5955; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25039.4]
  wire [1:0] _T_5956; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25040.4]
  wire [1:0] _T_5957; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25041.4]
  wire  _T_5958; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25042.4]
  wire  _T_5959; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25044.4]
  wire  _T_5961; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25046.4]
  wire  _T_5963; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25048.4]
  wire  _T_5964; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25049.4]
  wire  _T_5965; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25054.4]
  wire  _T_5966; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25055.4]
  wire  _T_5967; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25056.4]
  wire  _T_5969; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25058.4]
  wire  _T_5970; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25059.4]
  wire  _T_5981; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25076.4]
  wire  _T_5982; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25077.4]
  wire  _T_5984; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25079.4]
  wire  _T_5986; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25081.4]
  wire [1:0] _T_5987; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25082.4]
  wire [1:0] _T_5988; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25083.4]
  wire  _T_5989; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25084.4]
  wire  _T_5990; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25086.4]
  wire  _T_5992; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25088.4]
  wire  _T_5994; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25090.4]
  wire  _T_5995; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25091.4]
  wire  _T_5996; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25096.4]
  wire  _T_5997; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25097.4]
  wire  _T_5998; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25098.4]
  wire  _T_6000; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25100.4]
  wire  _T_6001; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25101.4]
  wire  _T_6012; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25118.4]
  wire  _T_6013; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25119.4]
  wire  _T_6015; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25121.4]
  wire  _T_6017; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25123.4]
  wire [1:0] _T_6018; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25124.4]
  wire [1:0] _T_6019; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25125.4]
  wire  _T_6020; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25126.4]
  wire  _T_6021; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25128.4]
  wire  _T_6023; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25130.4]
  wire  _T_6025; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25132.4]
  wire  _T_6026; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25133.4]
  wire  _T_6027; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25138.4]
  wire  _T_6028; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25139.4]
  wire  _T_6029; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25140.4]
  wire  _T_6031; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25142.4]
  wire  _T_6032; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25143.4]
  wire  _T_6043; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25160.4]
  wire  _T_6044; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25161.4]
  wire  _T_6046; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25163.4]
  wire  _T_6048; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25165.4]
  wire [1:0] _T_6049; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25166.4]
  wire [1:0] _T_6050; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25167.4]
  wire  _T_6051; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25168.4]
  wire  _T_6052; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25170.4]
  wire  _T_6054; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25172.4]
  wire  _T_6056; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25174.4]
  wire  _T_6057; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25175.4]
  wire  _T_6058; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25180.4]
  wire  _T_6059; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25181.4]
  wire  _T_6060; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25182.4]
  wire  _T_6062; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25184.4]
  wire  _T_6063; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25185.4]
  wire  _T_6074; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25202.4]
  wire  _T_6075; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25203.4]
  wire  _T_6077; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25205.4]
  wire  _T_6079; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25207.4]
  wire [1:0] _T_6080; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25208.4]
  wire [1:0] _T_6081; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25209.4]
  wire  _T_6082; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25210.4]
  wire  _T_6083; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25212.4]
  wire  _T_6085; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25214.4]
  wire  _T_6087; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25216.4]
  wire  _T_6088; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25217.4]
  wire  _T_6089; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25222.4]
  wire  _T_6090; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25223.4]
  wire  _T_6091; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25224.4]
  wire  _T_6093; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25226.4]
  wire  _T_6094; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25227.4]
  wire  _T_6105; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25244.4]
  wire  _T_6106; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25245.4]
  wire  _T_6108; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25247.4]
  wire  _T_6110; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25249.4]
  wire [1:0] _T_6111; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25250.4]
  wire [1:0] _T_6112; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25251.4]
  wire  _T_6113; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25252.4]
  wire  _T_6114; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25254.4]
  wire  _T_6116; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25256.4]
  wire  _T_6118; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25258.4]
  wire  _T_6119; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25259.4]
  wire  _T_6120; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25264.4]
  wire  _T_6121; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25265.4]
  wire  _T_6122; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25266.4]
  wire  _T_6124; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25268.4]
  wire  _T_6125; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25269.4]
  wire  _T_6136; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25286.4]
  wire  _T_6137; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25287.4]
  wire  _T_6139; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25289.4]
  wire  _T_6141; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25291.4]
  wire [1:0] _T_6142; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25292.4]
  wire [1:0] _T_6143; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25293.4]
  wire  _T_6144; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25294.4]
  wire  _T_6145; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25296.4]
  wire  _T_6147; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25298.4]
  wire  _T_6149; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25300.4]
  wire  _T_6150; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25301.4]
  wire  _T_6151; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25306.4]
  wire  _T_6152; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25307.4]
  wire  _T_6153; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25308.4]
  wire  _T_6155; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25310.4]
  wire  _T_6156; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25311.4]
  wire  _T_6167; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25328.4]
  wire  _T_6168; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25329.4]
  wire  _T_6170; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25331.4]
  wire  _T_6172; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25333.4]
  wire [1:0] _T_6173; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25334.4]
  wire [1:0] _T_6174; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25335.4]
  wire  _T_6175; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25336.4]
  wire  _T_6176; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25338.4]
  wire  _T_6178; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25340.4]
  wire  _T_6180; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25342.4]
  wire  _T_6181; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25343.4]
  wire  _T_6182; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25348.4]
  wire  _T_6183; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25349.4]
  wire  _T_6184; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25350.4]
  wire  _T_6186; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25352.4]
  wire  _T_6187; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25353.4]
  wire  _T_6198; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25370.4]
  wire  _T_6199; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25371.4]
  wire  _T_6201; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25373.4]
  wire  _T_6203; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25375.4]
  wire [1:0] _T_6204; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25376.4]
  wire [1:0] _T_6205; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25377.4]
  wire  _T_6206; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25378.4]
  wire  _T_6207; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25380.4]
  wire  _T_6209; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25382.4]
  wire  _T_6211; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25384.4]
  wire  _T_6212; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25385.4]
  wire  _T_6213; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25390.4]
  wire  _T_6214; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25391.4]
  wire  _T_6215; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25392.4]
  wire  _T_6217; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25394.4]
  wire  _T_6218; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25395.4]
  wire  _T_6229; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25412.4]
  wire  _T_6230; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25413.4]
  wire  _T_6232; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25415.4]
  wire  _T_6234; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25417.4]
  wire [1:0] _T_6235; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25418.4]
  wire [1:0] _T_6236; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25419.4]
  wire  _T_6237; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25420.4]
  wire  _T_6238; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25422.4]
  wire  _T_6240; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25424.4]
  wire  _T_6242; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25426.4]
  wire  _T_6243; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25427.4]
  wire  _T_6244; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25432.4]
  wire  _T_6245; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25433.4]
  wire  _T_6246; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25434.4]
  wire  _T_6248; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25436.4]
  wire  _T_6249; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25437.4]
  wire  _T_6260; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25454.4]
  wire  _T_6261; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25455.4]
  wire  _T_6263; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25457.4]
  wire  _T_6265; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25459.4]
  wire [1:0] _T_6266; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25460.4]
  wire [1:0] _T_6267; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25461.4]
  wire  _T_6268; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25462.4]
  wire  _T_6269; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25464.4]
  wire  _T_6271; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25466.4]
  wire  _T_6273; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25468.4]
  wire  _T_6274; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25469.4]
  wire  _T_6275; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25474.4]
  wire  _T_6276; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25475.4]
  wire  _T_6277; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25476.4]
  wire  _T_6279; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25478.4]
  wire  _T_6280; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25479.4]
  wire  _T_6291; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25496.4]
  wire  _T_6292; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25497.4]
  wire  _T_6294; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25499.4]
  wire  _T_6296; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25501.4]
  wire [1:0] _T_6297; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25502.4]
  wire [1:0] _T_6298; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25503.4]
  wire  _T_6299; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25504.4]
  wire  _T_6300; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25506.4]
  wire  _T_6302; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25508.4]
  wire  _T_6304; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25510.4]
  wire  _T_6305; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25511.4]
  wire  _T_6306; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25516.4]
  wire  _T_6307; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25517.4]
  wire  _T_6308; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25518.4]
  wire  _T_6310; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25520.4]
  wire  _T_6311; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25521.4]
  wire  _T_6322; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25538.4]
  wire  _T_6323; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25539.4]
  wire  _T_6325; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25541.4]
  wire  _T_6327; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25543.4]
  wire [1:0] _T_6328; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25544.4]
  wire [1:0] _T_6329; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25545.4]
  wire  _T_6330; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25546.4]
  wire  _T_6331; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25548.4]
  wire  _T_6333; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25550.4]
  wire  _T_6335; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25552.4]
  wire  _T_6336; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25553.4]
  wire  _T_6337; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25558.4]
  wire  _T_6338; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25559.4]
  wire  _T_6339; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25560.4]
  wire  _T_6341; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25562.4]
  wire  _T_6342; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25563.4]
  wire  _T_6353; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25580.4]
  wire  _T_6354; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25581.4]
  wire  _T_6356; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25583.4]
  wire  _T_6358; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25585.4]
  wire [1:0] _T_6359; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25586.4]
  wire [1:0] _T_6360; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25587.4]
  wire  _T_6361; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25588.4]
  wire  _T_6362; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25590.4]
  wire  _T_6364; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25592.4]
  wire  _T_6366; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25594.4]
  wire  _T_6367; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25595.4]
  wire  _T_6368; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25600.4]
  wire  _T_6369; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25601.4]
  wire  _T_6370; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25602.4]
  wire  _T_6372; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25604.4]
  wire  _T_6373; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25605.4]
  wire  _T_6384; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25622.4]
  wire  _T_6385; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25623.4]
  wire  _T_6387; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25625.4]
  wire  _T_6389; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25627.4]
  wire [1:0] _T_6390; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25628.4]
  wire [1:0] _T_6391; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25629.4]
  wire  _T_6392; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25630.4]
  wire  _T_6393; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25632.4]
  wire  _T_6395; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25634.4]
  wire  _T_6397; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25636.4]
  wire  _T_6398; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25637.4]
  wire  _T_6399; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25642.4]
  wire  _T_6400; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25643.4]
  wire  _T_6401; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25644.4]
  wire  _T_6403; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25646.4]
  wire  _T_6404; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25647.4]
  wire  _T_6415; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25664.4]
  wire  _T_6416; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25665.4]
  wire  _T_6418; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25667.4]
  wire  _T_6420; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25669.4]
  wire [1:0] _T_6421; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25670.4]
  wire [1:0] _T_6422; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25671.4]
  wire  _T_6423; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25672.4]
  wire  _T_6424; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25674.4]
  wire  _T_6426; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25676.4]
  wire  _T_6428; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25678.4]
  wire  _T_6429; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25679.4]
  wire  _T_6430; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25684.4]
  wire  _T_6431; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25685.4]
  wire  _T_6432; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25686.4]
  wire  _T_6434; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25688.4]
  wire  _T_6435; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25689.4]
  wire  _T_6446; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25706.4]
  wire  _T_6447; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25707.4]
  wire  _T_6449; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25709.4]
  wire  _T_6451; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25711.4]
  wire [1:0] _T_6452; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25712.4]
  wire [1:0] _T_6453; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25713.4]
  wire  _T_6454; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25714.4]
  wire  _T_6455; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25716.4]
  wire  _T_6457; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25718.4]
  wire  _T_6459; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25720.4]
  wire  _T_6460; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25721.4]
  wire  _T_6461; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25726.4]
  wire  _T_6462; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25727.4]
  wire  _T_6463; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25728.4]
  wire  _T_6465; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25730.4]
  wire  _T_6466; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25731.4]
  wire  _T_6477; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25748.4]
  wire  _T_6478; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25749.4]
  wire  _T_6480; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25751.4]
  wire  _T_6482; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25753.4]
  wire [1:0] _T_6483; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25754.4]
  wire [1:0] _T_6484; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25755.4]
  wire  _T_6485; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25756.4]
  wire  _T_6486; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25758.4]
  wire  _T_6488; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25760.4]
  wire  _T_6490; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25762.4]
  wire  _T_6491; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25763.4]
  wire  _T_6492; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25768.4]
  wire  _T_6493; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25769.4]
  wire  _T_6494; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25770.4]
  wire  _T_6496; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25772.4]
  wire  _T_6497; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25773.4]
  wire  _T_6508; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25790.4]
  wire  _T_6509; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25791.4]
  wire  _T_6511; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25793.4]
  wire  _T_6513; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25795.4]
  wire [1:0] _T_6514; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25796.4]
  wire [1:0] _T_6515; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25797.4]
  wire  _T_6516; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25798.4]
  wire  _T_6517; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25800.4]
  wire  _T_6519; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25802.4]
  wire  _T_6521; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25804.4]
  wire  _T_6522; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25805.4]
  wire  _T_6523; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25810.4]
  wire  _T_6524; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25811.4]
  wire  _T_6525; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25812.4]
  wire  _T_6527; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25814.4]
  wire  _T_6528; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25815.4]
  wire  _T_6539; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25832.4]
  wire  _T_6540; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25833.4]
  wire  _T_6542; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25835.4]
  wire  _T_6544; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25837.4]
  wire [1:0] _T_6545; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25838.4]
  wire [1:0] _T_6546; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25839.4]
  wire  _T_6547; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25840.4]
  wire  _T_6548; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25842.4]
  wire  _T_6550; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25844.4]
  wire  _T_6552; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25846.4]
  wire  _T_6553; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25847.4]
  wire  _T_6554; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25852.4]
  wire  _T_6555; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25853.4]
  wire  _T_6556; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25854.4]
  wire  _T_6558; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25856.4]
  wire  _T_6559; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25857.4]
  wire  _T_6570; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25874.4]
  wire  _T_6571; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25875.4]
  wire  _T_6573; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25877.4]
  wire  _T_6575; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25879.4]
  wire [1:0] _T_6576; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25880.4]
  wire [1:0] _T_6577; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25881.4]
  wire  _T_6578; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25882.4]
  wire  _T_6579; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25884.4]
  wire  _T_6581; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25886.4]
  wire  _T_6583; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25888.4]
  wire  _T_6584; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25889.4]
  wire  _T_6585; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25894.4]
  wire  _T_6586; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25895.4]
  wire  _T_6587; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25896.4]
  wire  _T_6589; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25898.4]
  wire  _T_6590; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25899.4]
  wire  _T_6601; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25916.4]
  wire  _T_6602; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25917.4]
  wire  _T_6604; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25919.4]
  wire  _T_6606; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25921.4]
  wire [1:0] _T_6607; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25922.4]
  wire [1:0] _T_6608; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25923.4]
  wire  _T_6609; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25924.4]
  wire  _T_6610; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25926.4]
  wire  _T_6612; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25928.4]
  wire  _T_6614; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25930.4]
  wire  _T_6615; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25931.4]
  wire  _T_6616; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25936.4]
  wire  _T_6617; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25937.4]
  wire  _T_6618; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25938.4]
  wire  _T_6620; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25940.4]
  wire  _T_6621; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25941.4]
  wire  _T_6632; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25958.4]
  wire  _T_6633; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25959.4]
  wire  _T_6635; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25961.4]
  wire  _T_6637; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25963.4]
  wire [1:0] _T_6638; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25964.4]
  wire [1:0] _T_6639; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25965.4]
  wire  _T_6640; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25966.4]
  wire  _T_6641; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25968.4]
  wire  _T_6643; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25970.4]
  wire  _T_6645; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25972.4]
  wire  _T_6646; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25973.4]
  wire  _T_6647; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25978.4]
  wire  _T_6648; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25979.4]
  wire  _T_6649; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25980.4]
  wire  _T_6651; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25982.4]
  wire  _T_6652; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25983.4]
  wire  _T_6663; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26000.4]
  wire  _T_6664; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26001.4]
  wire  _T_6666; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26003.4]
  wire  _T_6668; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26005.4]
  wire [1:0] _T_6669; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26006.4]
  wire [1:0] _T_6670; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26007.4]
  wire  _T_6671; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26008.4]
  wire  _T_6672; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26010.4]
  wire  _T_6674; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26012.4]
  wire  _T_6676; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26014.4]
  wire  _T_6677; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26015.4]
  wire  _T_6678; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26020.4]
  wire  _T_6679; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26021.4]
  wire  _T_6680; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26022.4]
  wire  _T_6682; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26024.4]
  wire  _T_6683; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26025.4]
  wire  _T_6694; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26042.4]
  wire  _T_6695; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26043.4]
  wire  _T_6697; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26045.4]
  wire  _T_6699; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26047.4]
  wire [1:0] _T_6700; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26048.4]
  wire [1:0] _T_6701; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26049.4]
  wire  _T_6702; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26050.4]
  wire  _T_6703; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26052.4]
  wire  _T_6705; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26054.4]
  wire  _T_6707; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26056.4]
  wire  _T_6708; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26057.4]
  wire  _T_6709; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26062.4]
  wire  _T_6710; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26063.4]
  wire  _T_6711; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26064.4]
  wire  _T_6713; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26066.4]
  wire  _T_6714; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26067.4]
  wire  _T_6725; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26084.4]
  wire  _T_6726; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26085.4]
  wire  _T_6728; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26087.4]
  wire  _T_6730; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26089.4]
  wire [1:0] _T_6731; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26090.4]
  wire [1:0] _T_6732; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26091.4]
  wire  _T_6733; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26092.4]
  wire  _T_6734; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26094.4]
  wire  _T_6736; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26096.4]
  wire  _T_6738; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26098.4]
  wire  _T_6739; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26099.4]
  wire  _T_6740; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26104.4]
  wire  _T_6741; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26105.4]
  wire  _T_6742; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26106.4]
  wire  _T_6744; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26108.4]
  wire  _T_6745; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26109.4]
  wire  _T_6756; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26126.4]
  wire  _T_6757; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26127.4]
  wire  _T_6759; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26129.4]
  wire  _T_6761; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26131.4]
  wire [1:0] _T_6762; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26132.4]
  wire [1:0] _T_6763; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26133.4]
  wire  _T_6764; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26134.4]
  wire  _T_6765; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26136.4]
  wire  _T_6767; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26138.4]
  wire  _T_6769; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26140.4]
  wire  _T_6770; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26141.4]
  wire  _T_6771; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26146.4]
  wire  _T_6772; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26147.4]
  wire  _T_6773; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26148.4]
  wire  _T_6775; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26150.4]
  wire  _T_6776; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26151.4]
  wire  _T_6787; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26168.4]
  wire  _T_6788; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26169.4]
  wire  _T_6790; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26171.4]
  wire  _T_6792; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26173.4]
  wire [1:0] _T_6793; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26174.4]
  wire [1:0] _T_6794; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26175.4]
  wire  _T_6795; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26176.4]
  wire  _T_6796; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26178.4]
  wire  _T_6798; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26180.4]
  wire  _T_6800; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26182.4]
  wire  _T_6801; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26183.4]
  wire  _T_6802; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26188.4]
  wire  _T_6803; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26189.4]
  wire  _T_6804; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26190.4]
  wire  _T_6806; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26192.4]
  wire  _T_6807; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26193.4]
  wire  _T_6818; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26210.4]
  wire  _T_6819; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26211.4]
  wire  _T_6821; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26213.4]
  wire  _T_6823; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26215.4]
  wire [1:0] _T_6824; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26216.4]
  wire [1:0] _T_6825; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26217.4]
  wire  _T_6826; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26218.4]
  wire  _T_6827; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26220.4]
  wire  _T_6829; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26222.4]
  wire  _T_6831; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26224.4]
  wire  _T_6832; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26225.4]
  wire  _T_6833; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26230.4]
  wire  _T_6834; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26231.4]
  wire  _T_6835; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26232.4]
  wire  _T_6837; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26234.4]
  wire  _T_6838; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26235.4]
  wire  _T_6849; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26252.4]
  wire  _T_6850; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26253.4]
  wire  _T_6852; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26255.4]
  wire  _T_6854; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26257.4]
  wire [1:0] _T_6855; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26258.4]
  wire [1:0] _T_6856; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26259.4]
  wire  _T_6857; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26260.4]
  wire  _T_6858; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26262.4]
  wire  _T_6860; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26264.4]
  wire  _T_6862; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26266.4]
  wire  _T_6863; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26267.4]
  wire  _T_6864; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26272.4]
  wire  _T_6865; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26273.4]
  wire  _T_6866; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26274.4]
  wire  _T_6868; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26276.4]
  wire  _T_6869; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26277.4]
  wire  _T_6880; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26294.4]
  wire  _T_6881; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26295.4]
  wire  _T_6883; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26297.4]
  wire  _T_6885; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26299.4]
  wire [1:0] _T_6886; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26300.4]
  wire [1:0] _T_6887; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26301.4]
  wire  _T_6888; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26302.4]
  wire  _T_6889; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26304.4]
  wire  _T_6891; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26306.4]
  wire  _T_6893; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26308.4]
  wire  _T_6894; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26309.4]
  wire  _T_6895; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26314.4]
  wire  _T_6896; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26315.4]
  wire  _T_6897; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26316.4]
  wire  _T_6899; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26318.4]
  wire  _T_6900; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26319.4]
  wire  _T_6911; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26336.4]
  wire  _T_6912; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26337.4]
  wire  _T_6914; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26339.4]
  wire  _T_6916; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26341.4]
  wire [1:0] _T_6917; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26342.4]
  wire [1:0] _T_6918; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26343.4]
  wire  _T_6919; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26344.4]
  wire  _T_6920; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26346.4]
  wire  _T_6922; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26348.4]
  wire  _T_6924; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26350.4]
  wire  _T_6925; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26351.4]
  wire  _T_6926; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26356.4]
  wire  _T_6927; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26357.4]
  wire  _T_6928; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26358.4]
  wire  _T_6930; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26360.4]
  wire  _T_6931; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26361.4]
  wire  _T_6942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26378.4]
  wire  _T_6943; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26379.4]
  wire  _T_6945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26381.4]
  wire  _T_6947; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26383.4]
  wire [1:0] _T_6948; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26384.4]
  wire [1:0] _T_6949; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26385.4]
  wire  _T_6950; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26386.4]
  wire  _T_6951; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26388.4]
  wire  _T_6953; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26390.4]
  wire  _T_6955; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26392.4]
  wire  _T_6956; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26393.4]
  wire  _T_6957; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26398.4]
  wire  _T_6958; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26399.4]
  wire  _T_6959; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26400.4]
  wire  _T_6961; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26402.4]
  wire  _T_6962; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26403.4]
  wire  _T_6973; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26420.4]
  wire  _T_6974; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26421.4]
  wire  _T_6976; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26423.4]
  wire  _T_6978; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26425.4]
  wire [1:0] _T_6979; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26426.4]
  wire [1:0] _T_6980; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26427.4]
  wire  _T_6981; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26428.4]
  wire  _T_6982; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26430.4]
  wire  _T_6984; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26432.4]
  wire  _T_6986; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26434.4]
  wire  _T_6987; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26435.4]
  wire  _T_6988; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26440.4]
  wire  _T_6989; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26441.4]
  wire  _T_6990; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26442.4]
  wire  _T_6992; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26444.4]
  wire  _T_6993; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26445.4]
  wire  _T_7004; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26462.4]
  wire  _T_7005; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26463.4]
  wire  _T_7007; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26465.4]
  wire  _T_7009; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26467.4]
  wire [1:0] _T_7010; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26468.4]
  wire [1:0] _T_7011; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26469.4]
  wire  _T_7012; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26470.4]
  wire  _T_7013; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26472.4]
  wire  _T_7015; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26474.4]
  wire  _T_7017; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26476.4]
  wire  _T_7018; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26477.4]
  wire  _T_7019; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26482.4]
  wire  _T_7020; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26483.4]
  wire  _T_7021; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26484.4]
  wire  _T_7023; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26486.4]
  wire  _T_7024; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26487.4]
  wire  _T_7035; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26504.4]
  wire  _T_7036; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26505.4]
  wire  _T_7038; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26507.4]
  wire  _T_7040; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26509.4]
  wire [1:0] _T_7041; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26510.4]
  wire [1:0] _T_7042; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26511.4]
  wire  _T_7043; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26512.4]
  wire  _T_7044; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26514.4]
  wire  _T_7046; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26516.4]
  wire  _T_7048; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26518.4]
  wire  _T_7049; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26519.4]
  wire  _T_7050; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26524.4]
  wire  _T_7051; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26525.4]
  wire  _T_7052; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26526.4]
  wire  _T_7054; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26528.4]
  wire  _T_7055; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26529.4]
  wire  _T_7066; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26546.4]
  wire  _T_7067; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26547.4]
  wire  _T_7069; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26549.4]
  wire  _T_7071; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26551.4]
  wire [1:0] _T_7072; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26552.4]
  wire [1:0] _T_7073; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26553.4]
  wire  _T_7074; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26554.4]
  wire  _T_7075; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26556.4]
  wire  _T_7077; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26558.4]
  wire  _T_7079; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26560.4]
  wire  _T_7080; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26561.4]
  wire  _T_7081; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26566.4]
  wire  _T_7082; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26567.4]
  wire  _T_7083; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26568.4]
  wire  _T_7085; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26570.4]
  wire  _T_7086; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26571.4]
  wire  _T_7097; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26588.4]
  wire  _T_7098; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26589.4]
  wire  _T_7100; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26591.4]
  wire  _T_7102; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26593.4]
  wire [1:0] _T_7103; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26594.4]
  wire [1:0] _T_7104; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26595.4]
  wire  _T_7105; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26596.4]
  wire  _T_7106; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26598.4]
  wire  _T_7108; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26600.4]
  wire  _T_7110; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26602.4]
  wire  _T_7111; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26603.4]
  wire  _T_7112; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26608.4]
  wire  _T_7113; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26609.4]
  wire  _T_7114; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26610.4]
  wire  _T_7116; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26612.4]
  wire  _T_7117; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26613.4]
  wire  _T_7128; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26630.4]
  wire  _T_7129; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26631.4]
  wire  _T_7131; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26633.4]
  wire  _T_7133; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26635.4]
  wire [1:0] _T_7134; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26636.4]
  wire [1:0] _T_7135; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26637.4]
  wire  _T_7136; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26638.4]
  wire  _T_7137; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26640.4]
  wire  _T_7139; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26642.4]
  wire  _T_7141; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26644.4]
  wire  _T_7142; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26645.4]
  wire  _T_7143; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26650.4]
  wire  _T_7144; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26651.4]
  wire  _T_7145; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26652.4]
  wire  _T_7147; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26654.4]
  wire  _T_7148; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26655.4]
  wire  _T_7159; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26672.4]
  wire  _T_7160; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26673.4]
  wire  _T_7162; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26675.4]
  wire  _T_7164; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26677.4]
  wire [1:0] _T_7165; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26678.4]
  wire [1:0] _T_7166; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26679.4]
  wire  _T_7167; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26680.4]
  wire  _T_7168; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26682.4]
  wire  _T_7170; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26684.4]
  wire  _T_7172; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26686.4]
  wire  _T_7173; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26687.4]
  wire  _T_7174; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26692.4]
  wire  _T_7175; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26693.4]
  wire  _T_7176; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26694.4]
  wire  _T_7178; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26696.4]
  wire  _T_7179; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26697.4]
  wire  _T_7190; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26714.4]
  wire  _T_7191; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26715.4]
  wire  _T_7193; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26717.4]
  wire  _T_7195; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26719.4]
  wire [1:0] _T_7196; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26720.4]
  wire [1:0] _T_7197; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26721.4]
  wire  _T_7198; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26722.4]
  wire  _T_7199; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26724.4]
  wire  _T_7201; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26726.4]
  wire  _T_7203; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26728.4]
  wire  _T_7204; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26729.4]
  wire  _T_7205; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26734.4]
  wire  _T_7206; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26735.4]
  wire  _T_7207; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26736.4]
  wire  _T_7209; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26738.4]
  wire  _T_7210; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26739.4]
  wire  _T_7221; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26756.4]
  wire  _T_7222; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26757.4]
  wire  _T_7224; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26759.4]
  wire  _T_7226; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26761.4]
  wire [1:0] _T_7227; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26762.4]
  wire [1:0] _T_7228; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26763.4]
  wire  _T_7229; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26764.4]
  wire  _T_7230; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26766.4]
  wire  _T_7232; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26768.4]
  wire  _T_7234; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26770.4]
  wire  _T_7235; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26771.4]
  wire  _T_7236; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26776.4]
  wire  _T_7237; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26777.4]
  wire  _T_7238; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26778.4]
  wire  _T_7240; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26780.4]
  wire  _T_7241; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26781.4]
  wire  _T_7252; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26798.4]
  wire  _T_7253; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26799.4]
  wire  _T_7255; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26801.4]
  wire  _T_7257; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26803.4]
  wire [1:0] _T_7258; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26804.4]
  wire [1:0] _T_7259; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26805.4]
  wire  _T_7260; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26806.4]
  wire  _T_7261; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26808.4]
  wire  _T_7263; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26810.4]
  wire  _T_7265; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26812.4]
  wire  _T_7266; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26813.4]
  wire  _T_7267; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26818.4]
  wire  _T_7268; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26819.4]
  wire  _T_7269; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26820.4]
  wire  _T_7271; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26822.4]
  wire  _T_7272; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26823.4]
  wire  _T_7283; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26840.4]
  wire  _T_7284; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26841.4]
  wire  _T_7286; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26843.4]
  wire  _T_7288; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26845.4]
  wire [1:0] _T_7289; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26846.4]
  wire [1:0] _T_7290; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26847.4]
  wire  _T_7291; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26848.4]
  wire  _T_7292; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26850.4]
  wire  _T_7294; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26852.4]
  wire  _T_7296; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26854.4]
  wire  _T_7297; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26855.4]
  wire  _T_7298; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26860.4]
  wire  _T_7299; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26861.4]
  wire  _T_7300; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26862.4]
  wire  _T_7302; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26864.4]
  wire  _T_7303; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26865.4]
  wire  _T_7314; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26882.4]
  wire  _T_7315; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26883.4]
  wire  _T_7317; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26885.4]
  wire  _T_7319; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26887.4]
  wire [1:0] _T_7320; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26888.4]
  wire [1:0] _T_7321; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26889.4]
  wire  _T_7322; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26890.4]
  wire  _T_7323; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26892.4]
  wire  _T_7325; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26894.4]
  wire  _T_7327; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26896.4]
  wire  _T_7328; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26897.4]
  wire  _T_7329; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26902.4]
  wire  _T_7330; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26903.4]
  wire  _T_7331; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26904.4]
  wire  _T_7333; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26906.4]
  wire  _T_7334; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26907.4]
  wire  _T_7345; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26924.4]
  wire  _T_7346; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26925.4]
  wire  _T_7348; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26927.4]
  wire  _T_7350; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26929.4]
  wire [1:0] _T_7351; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26930.4]
  wire [1:0] _T_7352; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26931.4]
  wire  _T_7353; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26932.4]
  wire  _T_7354; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26934.4]
  wire  _T_7356; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26936.4]
  wire  _T_7358; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26938.4]
  wire  _T_7359; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26939.4]
  wire  _T_7360; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26944.4]
  wire  _T_7361; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26945.4]
  wire  _T_7362; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26946.4]
  wire  _T_7364; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26948.4]
  wire  _T_7365; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26949.4]
  wire  _T_7376; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26966.4]
  wire  _T_7377; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26967.4]
  wire  _T_7379; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26969.4]
  wire  _T_7381; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26971.4]
  wire [1:0] _T_7382; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26972.4]
  wire [1:0] _T_7383; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26973.4]
  wire  _T_7384; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26974.4]
  wire  _T_7385; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26976.4]
  wire  _T_7387; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26978.4]
  wire  _T_7389; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26980.4]
  wire  _T_7390; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26981.4]
  wire  _T_7391; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26986.4]
  wire  _T_7392; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26987.4]
  wire  _T_7393; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26988.4]
  wire  _T_7395; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26990.4]
  wire  _T_7396; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26991.4]
  wire  _T_7407; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27008.4]
  wire  _T_7408; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27009.4]
  wire  _T_7410; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27011.4]
  wire  _T_7412; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27013.4]
  wire [1:0] _T_7413; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27014.4]
  wire [1:0] _T_7414; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27015.4]
  wire  _T_7415; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27016.4]
  wire  _T_7416; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27018.4]
  wire  _T_7418; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27020.4]
  wire  _T_7420; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27022.4]
  wire  _T_7421; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27023.4]
  wire  _T_7422; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27028.4]
  wire  _T_7423; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27029.4]
  wire  _T_7424; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27030.4]
  wire  _T_7426; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27032.4]
  wire  _T_7427; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27033.4]
  wire  _T_7438; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27050.4]
  wire  _T_7439; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27051.4]
  wire  _T_7441; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27053.4]
  wire  _T_7443; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27055.4]
  wire [1:0] _T_7444; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27056.4]
  wire [1:0] _T_7445; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27057.4]
  wire  _T_7446; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27058.4]
  wire  _T_7447; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27060.4]
  wire  _T_7449; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27062.4]
  wire  _T_7451; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27064.4]
  wire  _T_7452; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27065.4]
  wire  _T_7453; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27070.4]
  wire  _T_7454; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27071.4]
  wire  _T_7455; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27072.4]
  wire  _T_7457; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27074.4]
  wire  _T_7458; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27075.4]
  wire  _T_7469; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27092.4]
  wire  _T_7470; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27093.4]
  wire  _T_7472; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27095.4]
  wire  _T_7474; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27097.4]
  wire [1:0] _T_7475; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27098.4]
  wire [1:0] _T_7476; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27099.4]
  wire  _T_7477; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27100.4]
  wire  _T_7478; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27102.4]
  wire  _T_7480; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27104.4]
  wire  _T_7482; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27106.4]
  wire  _T_7483; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27107.4]
  wire  _T_7484; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27112.4]
  wire  _T_7485; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27113.4]
  wire  _T_7486; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27114.4]
  wire  _T_7488; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27116.4]
  wire  _T_7489; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27117.4]
  wire  _T_7500; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27134.4]
  wire  _T_7501; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27135.4]
  wire  _T_7503; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27137.4]
  wire  _T_7505; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27139.4]
  wire [1:0] _T_7506; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27140.4]
  wire [1:0] _T_7507; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27141.4]
  wire  _T_7508; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27142.4]
  wire  _T_7509; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27144.4]
  wire  _T_7511; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27146.4]
  wire  _T_7513; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27148.4]
  wire  _T_7514; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27149.4]
  wire  _T_7515; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27154.4]
  wire  _T_7516; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27155.4]
  wire  _T_7517; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27156.4]
  wire  _T_7519; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27158.4]
  wire  _T_7520; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27159.4]
  wire  _T_7531; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27176.4]
  wire  _T_7532; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27177.4]
  wire  _T_7534; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27179.4]
  wire  _T_7536; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27181.4]
  wire [1:0] _T_7537; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27182.4]
  wire [1:0] _T_7538; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27183.4]
  wire  _T_7539; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27184.4]
  wire  _T_7540; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27186.4]
  wire  _T_7542; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27188.4]
  wire  _T_7544; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27190.4]
  wire  _T_7545; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27191.4]
  wire  _T_7546; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27196.4]
  wire  _T_7547; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27197.4]
  wire  _T_7548; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27198.4]
  wire  _T_7550; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27200.4]
  wire  _T_7551; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27201.4]
  wire  _T_7562; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27218.4]
  wire  _T_7563; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27219.4]
  wire  _T_7565; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27221.4]
  wire  _T_7567; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27223.4]
  wire [1:0] _T_7568; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27224.4]
  wire [1:0] _T_7569; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27225.4]
  wire  _T_7570; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27226.4]
  wire  _T_7571; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27228.4]
  wire  _T_7573; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27230.4]
  wire  _T_7575; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27232.4]
  wire  _T_7576; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27233.4]
  wire  _T_7577; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27238.4]
  wire  _T_7578; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27239.4]
  wire  _T_7579; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27240.4]
  wire  _T_7581; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27242.4]
  wire  _T_7582; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27243.4]
  wire  _T_7593; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27260.4]
  wire  _T_7594; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27261.4]
  wire  _T_7596; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27263.4]
  wire  _T_7598; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27265.4]
  wire [1:0] _T_7599; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27266.4]
  wire [1:0] _T_7600; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27267.4]
  wire  _T_7601; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27268.4]
  wire  _T_7602; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27270.4]
  wire  _T_7604; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27272.4]
  wire  _T_7606; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27274.4]
  wire  _T_7607; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27275.4]
  wire  _T_7608; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27280.4]
  wire  _T_7609; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27281.4]
  wire  _T_7610; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27282.4]
  wire  _T_7612; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27284.4]
  wire  _T_7613; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27285.4]
  wire  _T_7624; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27302.4]
  wire  _T_7625; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27303.4]
  wire  _T_7627; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27305.4]
  wire  _T_7629; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27307.4]
  wire [1:0] _T_7630; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27308.4]
  wire [1:0] _T_7631; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27309.4]
  wire  _T_7632; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27310.4]
  wire  _T_7633; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27312.4]
  wire  _T_7635; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27314.4]
  wire  _T_7637; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27316.4]
  wire  _T_7638; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27317.4]
  wire  _T_7639; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27322.4]
  wire  _T_7640; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27323.4]
  wire  _T_7641; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27324.4]
  wire  _T_7643; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27326.4]
  wire  _T_7644; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27327.4]
  wire  _T_7655; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27344.4]
  wire  _T_7656; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27345.4]
  wire  _T_7658; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27347.4]
  wire  _T_7660; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27349.4]
  wire [1:0] _T_7661; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27350.4]
  wire [1:0] _T_7662; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27351.4]
  wire  _T_7663; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27352.4]
  wire  _T_7664; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27354.4]
  wire  _T_7666; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27356.4]
  wire  _T_7668; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27358.4]
  wire  _T_7669; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27359.4]
  wire  _T_7670; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27364.4]
  wire  _T_7671; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27365.4]
  wire  _T_7672; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27366.4]
  wire  _T_7674; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27368.4]
  wire  _T_7675; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27369.4]
  wire  _T_7686; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27386.4]
  wire  _T_7687; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27387.4]
  wire  _T_7689; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27389.4]
  wire  _T_7691; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27391.4]
  wire [1:0] _T_7692; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27392.4]
  wire [1:0] _T_7693; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27393.4]
  wire  _T_7694; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27394.4]
  wire  _T_7695; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27396.4]
  wire  _T_7697; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27398.4]
  wire  _T_7699; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27400.4]
  wire  _T_7700; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27401.4]
  wire  _T_7701; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27406.4]
  wire  _T_7702; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27407.4]
  wire  _T_7703; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27408.4]
  wire  _T_7705; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27410.4]
  wire  _T_7706; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27411.4]
  wire  _T_7717; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27428.4]
  wire  _T_7718; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27429.4]
  wire  _T_7720; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27431.4]
  wire  _T_7722; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27433.4]
  wire [1:0] _T_7723; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27434.4]
  wire [1:0] _T_7724; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27435.4]
  wire  _T_7725; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27436.4]
  wire  _T_7726; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27438.4]
  wire  _T_7728; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27440.4]
  wire  _T_7730; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27442.4]
  wire  _T_7731; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27443.4]
  wire  _T_7732; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27448.4]
  wire  _T_7733; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27449.4]
  wire  _T_7734; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27450.4]
  wire  _T_7736; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27452.4]
  wire  _T_7737; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27453.4]
  wire  _T_7748; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27470.4]
  wire  _T_7749; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27471.4]
  wire  _T_7751; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27473.4]
  wire  _T_7753; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27475.4]
  wire [1:0] _T_7754; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27476.4]
  wire [1:0] _T_7755; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27477.4]
  wire  _T_7756; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27478.4]
  wire  _T_7757; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27480.4]
  wire  _T_7759; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27482.4]
  wire  _T_7761; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27484.4]
  wire  _T_7762; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27485.4]
  wire  _T_7763; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27490.4]
  wire  _T_7764; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27491.4]
  wire  _T_7765; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27492.4]
  wire  _T_7767; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27494.4]
  wire  _T_7768; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27495.4]
  wire  _T_7779; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27512.4]
  wire  _T_7780; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27513.4]
  wire  _T_7782; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27515.4]
  wire  _T_7784; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27517.4]
  wire [1:0] _T_7785; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27518.4]
  wire [1:0] _T_7786; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27519.4]
  wire  _T_7787; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27520.4]
  wire  _T_7788; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27522.4]
  wire  _T_7790; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27524.4]
  wire  _T_7792; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27526.4]
  wire  _T_7793; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27527.4]
  wire  _T_7794; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27532.4]
  wire  _T_7795; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27533.4]
  wire  _T_7796; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27534.4]
  wire  _T_7798; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27536.4]
  wire  _T_7799; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27537.4]
  wire  _T_7810; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27554.4]
  wire  _T_7811; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27555.4]
  wire  _T_7813; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27557.4]
  wire  _T_7815; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27559.4]
  wire [1:0] _T_7816; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27560.4]
  wire [1:0] _T_7817; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27561.4]
  wire  _T_7818; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27562.4]
  wire  _T_7819; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27564.4]
  wire  _T_7821; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27566.4]
  wire  _T_7823; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27568.4]
  wire  _T_7824; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27569.4]
  wire  _T_7825; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27574.4]
  wire  _T_7826; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27575.4]
  wire  _T_7827; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27576.4]
  wire  _T_7829; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27578.4]
  wire  _T_7830; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27579.4]
  wire  _T_7841; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27596.4]
  wire  _T_7842; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27597.4]
  wire  _T_7844; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27599.4]
  wire  _T_7846; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27601.4]
  wire [1:0] _T_7847; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27602.4]
  wire [1:0] _T_7848; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27603.4]
  wire  _T_7849; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27604.4]
  wire  _T_7850; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27606.4]
  wire  _T_7852; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27608.4]
  wire  _T_7854; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27610.4]
  wire  _T_7855; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27611.4]
  wire  _T_7856; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27616.4]
  wire  _T_7857; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27617.4]
  wire  _T_7858; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27618.4]
  wire  _T_7860; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27620.4]
  wire  _T_7861; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27621.4]
  wire  _T_7872; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27638.4]
  wire  _T_7873; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27639.4]
  wire  _T_7875; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27641.4]
  wire  _T_7877; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27643.4]
  wire [1:0] _T_7878; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27644.4]
  wire [1:0] _T_7879; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27645.4]
  wire  _T_7880; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27646.4]
  wire  _T_7881; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27648.4]
  wire  _T_7883; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27650.4]
  wire  _T_7885; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27652.4]
  wire  _T_7886; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27653.4]
  wire  _T_7887; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27658.4]
  wire  _T_7888; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27659.4]
  wire  _T_7889; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27660.4]
  wire  _T_7891; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27662.4]
  wire  _T_7892; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27663.4]
  wire  _T_7903; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27680.4]
  wire  _T_7904; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27681.4]
  wire  _T_7906; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27683.4]
  wire  _T_7908; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27685.4]
  wire [1:0] _T_7909; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27686.4]
  wire [1:0] _T_7910; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27687.4]
  wire  _T_7911; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27688.4]
  wire  _T_7912; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27690.4]
  wire  _T_7914; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27692.4]
  wire  _T_7916; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27694.4]
  wire  _T_7917; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27695.4]
  wire  _T_7918; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27700.4]
  wire  _T_7919; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27701.4]
  wire  _T_7920; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27702.4]
  wire  _T_7922; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27704.4]
  wire  _T_7923; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27705.4]
  wire  _T_7934; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27722.4]
  wire  _T_7935; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27723.4]
  wire  _T_7937; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27725.4]
  wire  _T_7939; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27727.4]
  wire [1:0] _T_7940; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27728.4]
  wire [1:0] _T_7941; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27729.4]
  wire  _T_7942; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27730.4]
  wire  _T_7943; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27732.4]
  wire  _T_7945; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27734.4]
  wire  _T_7947; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27736.4]
  wire  _T_7948; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27737.4]
  wire  _T_7949; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27742.4]
  wire  _T_7950; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27743.4]
  wire  _T_7951; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27744.4]
  wire  _T_7953; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27746.4]
  wire  _T_7954; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27747.4]
  wire  _T_7965; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27764.4]
  wire  _T_7966; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27765.4]
  wire  _T_7968; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27767.4]
  wire  _T_7970; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27769.4]
  wire [1:0] _T_7971; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27770.4]
  wire [1:0] _T_7972; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27771.4]
  wire  _T_7973; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27772.4]
  wire  _T_7974; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27774.4]
  wire  _T_7976; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27776.4]
  wire  _T_7978; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27778.4]
  wire  _T_7979; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27779.4]
  wire  _T_7980; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27784.4]
  wire  _T_7981; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27785.4]
  wire  _T_7982; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27786.4]
  wire  _T_7984; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27788.4]
  wire  _T_7985; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27789.4]
  wire  _T_7996; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27806.4]
  wire  _T_7997; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27807.4]
  wire  _T_7999; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27809.4]
  wire  _T_8001; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27811.4]
  wire [1:0] _T_8002; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27812.4]
  wire [1:0] _T_8003; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27813.4]
  wire  _T_8004; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27814.4]
  wire  _T_8005; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27816.4]
  wire  _T_8007; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27818.4]
  wire  _T_8009; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27820.4]
  wire  _T_8010; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27821.4]
  wire  _T_8011; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27826.4]
  wire  _T_8012; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27827.4]
  wire  _T_8013; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27828.4]
  wire  _T_8015; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27830.4]
  wire  _T_8016; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27831.4]
  wire  _T_8027; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27848.4]
  wire  _T_8028; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27849.4]
  wire  _T_8030; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27851.4]
  wire  _T_8032; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27853.4]
  wire [1:0] _T_8033; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27854.4]
  wire [1:0] _T_8034; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27855.4]
  wire  _T_8035; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27856.4]
  wire  _T_8036; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27858.4]
  wire  _T_8038; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27860.4]
  wire  _T_8040; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27862.4]
  wire  _T_8041; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27863.4]
  wire  _T_8042; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27868.4]
  wire  _T_8043; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27869.4]
  wire  _T_8044; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27870.4]
  wire  _T_8046; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27872.4]
  wire  _T_8047; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27873.4]
  wire  _T_8058; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27890.4]
  wire  _T_8059; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27891.4]
  wire  _T_8061; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27893.4]
  wire  _T_8063; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27895.4]
  wire [1:0] _T_8064; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27896.4]
  wire [1:0] _T_8065; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27897.4]
  wire  _T_8066; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27898.4]
  wire  _T_8067; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27900.4]
  wire  _T_8069; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27902.4]
  wire  _T_8071; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27904.4]
  wire  _T_8072; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27905.4]
  wire  _T_8073; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27910.4]
  wire  _T_8074; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27911.4]
  wire  _T_8075; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27912.4]
  wire  _T_8077; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27914.4]
  wire  _T_8078; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27915.4]
  wire  _T_8089; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27932.4]
  wire  _T_8090; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27933.4]
  wire  _T_8092; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27935.4]
  wire  _T_8094; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27937.4]
  wire [1:0] _T_8095; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27938.4]
  wire [1:0] _T_8096; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27939.4]
  wire  _T_8097; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27940.4]
  wire  _T_8098; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27942.4]
  wire  _T_8100; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27944.4]
  wire  _T_8102; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27946.4]
  wire  _T_8103; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27947.4]
  wire  _T_8104; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27952.4]
  wire  _T_8105; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27953.4]
  wire  _T_8106; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27954.4]
  wire  _T_8108; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27956.4]
  wire  _T_8109; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27957.4]
  wire  _T_8120; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27974.4]
  wire  _T_8121; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27975.4]
  wire  _T_8123; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27977.4]
  wire  _T_8125; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27979.4]
  wire [1:0] _T_8126; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27980.4]
  wire [1:0] _T_8127; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27981.4]
  wire  _T_8128; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27982.4]
  wire  _T_8129; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27984.4]
  wire  _T_8131; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27986.4]
  wire  _T_8133; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27988.4]
  wire  _T_8134; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27989.4]
  wire  _T_8135; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27994.4]
  wire  _T_8136; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27995.4]
  wire  _T_8137; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27996.4]
  wire  _T_8139; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27998.4]
  wire  _T_8140; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27999.4]
  wire  _T_8151; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28016.4]
  wire  _T_8152; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28017.4]
  wire  _T_8154; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28019.4]
  wire  _T_8156; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28021.4]
  wire [1:0] _T_8157; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28022.4]
  wire [1:0] _T_8158; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28023.4]
  wire  _T_8159; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28024.4]
  wire  _T_8160; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28026.4]
  wire  _T_8162; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28028.4]
  wire  _T_8164; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28030.4]
  wire  _T_8165; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28031.4]
  wire  _T_8166; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28036.4]
  wire  _T_8167; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28037.4]
  wire  _T_8168; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28038.4]
  wire  _T_8170; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28040.4]
  wire  _T_8171; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28041.4]
  wire  _T_8182; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28058.4]
  wire  _T_8183; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28059.4]
  wire  _T_8185; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28061.4]
  wire  _T_8187; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28063.4]
  wire [1:0] _T_8188; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28064.4]
  wire [1:0] _T_8189; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28065.4]
  wire  _T_8190; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28066.4]
  wire  _T_8191; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28068.4]
  wire  _T_8193; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28070.4]
  wire  _T_8195; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28072.4]
  wire  _T_8196; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28073.4]
  wire  _T_8197; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28078.4]
  wire  _T_8198; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28079.4]
  wire  _T_8199; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28080.4]
  wire  _T_8201; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28082.4]
  wire  _T_8202; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28083.4]
  wire  _T_8213; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28100.4]
  wire  _T_8214; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28101.4]
  wire  _T_8216; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28103.4]
  wire  _T_8218; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28105.4]
  wire [1:0] _T_8219; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28106.4]
  wire [1:0] _T_8220; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28107.4]
  wire  _T_8221; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28108.4]
  wire  _T_8222; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28110.4]
  wire  _T_8224; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28112.4]
  wire  _T_8226; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28114.4]
  wire  _T_8227; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28115.4]
  wire  _T_8228; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28120.4]
  wire  _T_8229; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28121.4]
  wire  _T_8230; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28122.4]
  wire  _T_8232; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28124.4]
  wire  _T_8233; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28125.4]
  wire  _T_8244; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28142.4]
  wire  _T_8245; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28143.4]
  wire  _T_8247; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28145.4]
  wire  _T_8249; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28147.4]
  wire [1:0] _T_8250; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28148.4]
  wire [1:0] _T_8251; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28149.4]
  wire  _T_8252; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28150.4]
  wire  _T_8253; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28152.4]
  wire  _T_8255; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28154.4]
  wire  _T_8257; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28156.4]
  wire  _T_8258; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28157.4]
  wire  _T_8259; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28162.4]
  wire  _T_8260; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28163.4]
  wire  _T_8261; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28164.4]
  wire  _T_8263; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28166.4]
  wire  _T_8264; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28167.4]
  wire  _T_8275; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28184.4]
  wire  _T_8276; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28185.4]
  wire  _T_8278; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28187.4]
  wire  _T_8280; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28189.4]
  wire [1:0] _T_8281; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28190.4]
  wire [1:0] _T_8282; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28191.4]
  wire  _T_8283; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28192.4]
  wire  _T_8284; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28194.4]
  wire  _T_8286; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28196.4]
  wire  _T_8288; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28198.4]
  wire  _T_8289; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28199.4]
  wire  _T_8290; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28204.4]
  wire  _T_8291; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28205.4]
  wire  _T_8292; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28206.4]
  wire  _T_8294; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28208.4]
  wire  _T_8295; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28209.4]
  wire  _T_8306; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28226.4]
  wire  _T_8307; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28227.4]
  wire  _T_8309; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28229.4]
  wire  _T_8311; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28231.4]
  wire [1:0] _T_8312; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28232.4]
  wire [1:0] _T_8313; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28233.4]
  wire  _T_8314; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28234.4]
  wire  _T_8315; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28236.4]
  wire  _T_8317; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28238.4]
  wire  _T_8319; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28240.4]
  wire  _T_8320; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28241.4]
  wire  _T_8321; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28246.4]
  wire  _T_8322; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28247.4]
  wire  _T_8323; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28248.4]
  wire  _T_8325; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28250.4]
  wire  _T_8326; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28251.4]
  wire  _T_8337; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28268.4]
  wire  _T_8338; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28269.4]
  wire  _T_8340; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28271.4]
  wire  _T_8342; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28273.4]
  wire [1:0] _T_8343; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28274.4]
  wire [1:0] _T_8344; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28275.4]
  wire  _T_8345; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28276.4]
  wire  _T_8346; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28278.4]
  wire  _T_8348; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28280.4]
  wire  _T_8350; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28282.4]
  wire  _T_8351; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28283.4]
  wire  _T_8352; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28288.4]
  wire  _T_8353; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28289.4]
  wire  _T_8354; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28290.4]
  wire  _T_8356; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28292.4]
  wire  _T_8357; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28293.4]
  wire  _T_8368; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28310.4]
  wire  _T_8369; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28311.4]
  wire  _T_8371; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28313.4]
  wire  _T_8373; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28315.4]
  wire [1:0] _T_8374; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28316.4]
  wire [1:0] _T_8375; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28317.4]
  wire  _T_8376; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28318.4]
  wire  _T_8377; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28320.4]
  wire  _T_8379; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28322.4]
  wire  _T_8381; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28324.4]
  wire  _T_8382; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28325.4]
  wire  _T_8383; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28330.4]
  wire  _T_8384; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28331.4]
  wire  _T_8385; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28332.4]
  wire  _T_8387; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28334.4]
  wire  _T_8388; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28335.4]
  wire  _T_8399; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28352.4]
  wire  _T_8400; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28353.4]
  wire  _T_8402; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28355.4]
  wire  _T_8404; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28357.4]
  wire [1:0] _T_8405; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28358.4]
  wire [1:0] _T_8406; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28359.4]
  wire  _T_8407; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28360.4]
  wire  _T_8408; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28362.4]
  wire  _T_8410; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28364.4]
  wire  _T_8412; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28366.4]
  wire  _T_8413; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28367.4]
  wire  _T_8414; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28372.4]
  wire  _T_8415; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28373.4]
  wire  _T_8416; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28374.4]
  wire  _T_8418; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28376.4]
  wire  _T_8419; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28377.4]
  wire  _T_8430; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28394.4]
  wire  _T_8431; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28395.4]
  wire  _T_8433; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28397.4]
  wire  _T_8435; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28399.4]
  wire [1:0] _T_8436; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28400.4]
  wire [1:0] _T_8437; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28401.4]
  wire  _T_8438; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28402.4]
  wire  _T_8439; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28404.4]
  wire  _T_8441; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28406.4]
  wire  _T_8443; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28408.4]
  wire  _T_8444; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28409.4]
  wire  _T_8445; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28414.4]
  wire  _T_8446; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28415.4]
  wire  _T_8447; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28416.4]
  wire  _T_8449; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28418.4]
  wire  _T_8450; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28419.4]
  wire  _T_8461; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28436.4]
  wire  _T_8462; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28437.4]
  wire  _T_8464; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28439.4]
  wire  _T_8466; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28441.4]
  wire [1:0] _T_8467; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28442.4]
  wire [1:0] _T_8468; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28443.4]
  wire  _T_8469; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28444.4]
  wire  _T_8470; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28446.4]
  wire  _T_8472; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28448.4]
  wire  _T_8474; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28450.4]
  wire  _T_8475; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28451.4]
  wire  _T_8476; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28456.4]
  wire  _T_8477; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28457.4]
  wire  _T_8478; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28458.4]
  wire  _T_8480; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28460.4]
  wire  _T_8481; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28461.4]
  wire  _T_8492; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28478.4]
  wire  _T_8493; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28479.4]
  wire  _T_8495; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28481.4]
  wire  _T_8497; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28483.4]
  wire [1:0] _T_8498; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28484.4]
  wire [1:0] _T_8499; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28485.4]
  wire  _T_8500; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28486.4]
  wire  _T_8501; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28488.4]
  wire  _T_8503; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28490.4]
  wire  _T_8505; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28492.4]
  wire  _T_8506; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28493.4]
  wire  _T_8507; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28498.4]
  wire  _T_8508; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28499.4]
  wire  _T_8509; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28500.4]
  wire  _T_8511; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28502.4]
  wire  _T_8512; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28503.4]
  wire  _T_8523; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28520.4]
  wire  _T_8524; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28521.4]
  wire  _T_8526; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28523.4]
  wire  _T_8528; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28525.4]
  wire [1:0] _T_8529; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28526.4]
  wire [1:0] _T_8530; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28527.4]
  wire  _T_8531; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28528.4]
  wire  _T_8532; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28530.4]
  wire  _T_8534; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28532.4]
  wire  _T_8536; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28534.4]
  wire  _T_8537; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28535.4]
  wire  _T_8538; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28540.4]
  wire  _T_8539; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28541.4]
  wire  _T_8540; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28542.4]
  wire  _T_8542; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28544.4]
  wire  _T_8543; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28545.4]
  wire  _T_8554; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28562.4]
  wire  _T_8555; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28563.4]
  wire  _T_8557; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28565.4]
  wire  _T_8559; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28567.4]
  wire [1:0] _T_8560; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28568.4]
  wire [1:0] _T_8561; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28569.4]
  wire  _T_8562; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28570.4]
  wire  _T_8563; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28572.4]
  wire  _T_8565; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28574.4]
  wire  _T_8567; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28576.4]
  wire  _T_8568; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28577.4]
  wire  _T_8569; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28582.4]
  wire  _T_8570; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28583.4]
  wire  _T_8571; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28584.4]
  wire  _T_8573; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28586.4]
  wire  _T_8574; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28587.4]
  wire  _T_8585; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28604.4]
  wire  _T_8586; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28605.4]
  wire  _T_8588; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28607.4]
  wire  _T_8590; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28609.4]
  wire [1:0] _T_8591; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28610.4]
  wire [1:0] _T_8592; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28611.4]
  wire  _T_8593; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28612.4]
  wire  _T_8594; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28614.4]
  wire  _T_8596; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28616.4]
  wire  _T_8598; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28618.4]
  wire  _T_8599; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28619.4]
  wire  _T_8600; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28624.4]
  wire  _T_8601; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28625.4]
  wire  _T_8602; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28626.4]
  wire  _T_8604; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28628.4]
  wire  _T_8605; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28629.4]
  wire  _T_8616; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28646.4]
  wire  _T_8617; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28647.4]
  wire  _T_8619; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28649.4]
  wire  _T_8621; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28651.4]
  wire [1:0] _T_8622; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28652.4]
  wire [1:0] _T_8623; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28653.4]
  wire  _T_8624; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28654.4]
  wire  _T_8625; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28656.4]
  wire  _T_8627; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28658.4]
  wire  _T_8629; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28660.4]
  wire  _T_8630; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28661.4]
  wire  _T_8631; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28666.4]
  wire  _T_8632; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28667.4]
  wire  _T_8633; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28668.4]
  wire  _T_8635; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28670.4]
  wire  _T_8636; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28671.4]
  wire  _T_8647; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28688.4]
  wire  _T_8648; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28689.4]
  wire  _T_8650; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28691.4]
  wire  _T_8652; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28693.4]
  wire [1:0] _T_8653; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28694.4]
  wire [1:0] _T_8654; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28695.4]
  wire  _T_8655; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28696.4]
  wire  _T_8656; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28698.4]
  wire  _T_8658; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28700.4]
  wire  _T_8660; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28702.4]
  wire  _T_8661; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28703.4]
  wire  _T_8662; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28708.4]
  wire  _T_8663; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28709.4]
  wire  _T_8664; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28710.4]
  wire  _T_8666; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28712.4]
  wire  _T_8667; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28713.4]
  wire  _T_8678; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28730.4]
  wire  _T_8679; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28731.4]
  wire  _T_8681; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28733.4]
  wire  _T_8683; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28735.4]
  wire [1:0] _T_8684; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28736.4]
  wire [1:0] _T_8685; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28737.4]
  wire  _T_8686; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28738.4]
  wire  _T_8687; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28740.4]
  wire  _T_8689; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28742.4]
  wire  _T_8691; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28744.4]
  wire  _T_8692; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28745.4]
  wire  _T_8693; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28750.4]
  wire  _T_8694; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28751.4]
  wire  _T_8695; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28752.4]
  wire  _T_8697; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28754.4]
  wire  _T_8698; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28755.4]
  wire  _T_8709; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28772.4]
  wire  _T_8710; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28773.4]
  wire  _T_8712; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28775.4]
  wire  _T_8714; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28777.4]
  wire [1:0] _T_8715; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28778.4]
  wire [1:0] _T_8716; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28779.4]
  wire  _T_8717; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28780.4]
  wire  _T_8718; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28782.4]
  wire  _T_8720; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28784.4]
  wire  _T_8722; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28786.4]
  wire  _T_8723; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28787.4]
  wire  _T_8724; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28792.4]
  wire  _T_8725; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28793.4]
  wire  _T_8726; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28794.4]
  wire  _T_8728; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28796.4]
  wire  _T_8729; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28797.4]
  wire  _T_8740; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28814.4]
  wire  _T_8741; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28815.4]
  wire  _T_8743; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28817.4]
  wire  _T_8745; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28819.4]
  wire [1:0] _T_8746; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28820.4]
  wire [1:0] _T_8747; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28821.4]
  wire  _T_8748; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28822.4]
  wire  _T_8749; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28824.4]
  wire  _T_8751; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28826.4]
  wire  _T_8753; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28828.4]
  wire  _T_8754; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28829.4]
  wire  _T_8755; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28834.4]
  wire  _T_8756; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28835.4]
  wire  _T_8757; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28836.4]
  wire  _T_8759; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28838.4]
  wire  _T_8760; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28839.4]
  wire  _T_8771; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28856.4]
  wire  _T_8772; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28857.4]
  wire  _T_8774; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28859.4]
  wire  _T_8776; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28861.4]
  wire [1:0] _T_8777; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28862.4]
  wire [1:0] _T_8778; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28863.4]
  wire  _T_8779; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28864.4]
  wire  _T_8780; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28866.4]
  wire  _T_8782; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28868.4]
  wire  _T_8784; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28870.4]
  wire  _T_8785; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28871.4]
  wire  _T_8786; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28876.4]
  wire  _T_8787; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28877.4]
  wire  _T_8788; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28878.4]
  wire  _T_8790; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28880.4]
  wire  _T_8791; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28881.4]
  wire  _T_8802; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28898.4]
  wire  _T_8803; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28899.4]
  wire  _T_8805; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28901.4]
  wire  _T_8807; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28903.4]
  wire [1:0] _T_8808; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28904.4]
  wire [1:0] _T_8809; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28905.4]
  wire  _T_8810; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28906.4]
  wire  _T_8811; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28908.4]
  wire  _T_8813; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28910.4]
  wire  _T_8815; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28912.4]
  wire  _T_8816; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28913.4]
  wire  _T_8817; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28918.4]
  wire  _T_8818; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28919.4]
  wire  _T_8819; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28920.4]
  wire  _T_8821; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28922.4]
  wire  _T_8822; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28923.4]
  wire  _T_8833; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28940.4]
  wire  _T_8834; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28941.4]
  wire  _T_8836; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28943.4]
  wire  _T_8838; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28945.4]
  wire [1:0] _T_8839; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28946.4]
  wire [1:0] _T_8840; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28947.4]
  wire  _T_8841; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28948.4]
  wire  _T_8842; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28950.4]
  wire  _T_8844; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28952.4]
  wire  _T_8846; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28954.4]
  wire  _T_8847; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28955.4]
  wire  _T_8848; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28960.4]
  wire  _T_8849; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28961.4]
  wire  _T_8850; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28962.4]
  wire  _T_8852; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28964.4]
  wire  _T_8853; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28965.4]
  wire  _T_8864; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28982.4]
  wire  _T_8865; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28983.4]
  wire  _T_8867; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28985.4]
  wire  _T_8869; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28987.4]
  wire [1:0] _T_8870; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28988.4]
  wire [1:0] _T_8871; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28989.4]
  wire  _T_8872; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28990.4]
  wire  _T_8873; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28992.4]
  wire  _T_8875; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28994.4]
  wire  _T_8877; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28996.4]
  wire  _T_8878; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28997.4]
  wire  _T_8879; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29002.4]
  wire  _T_8880; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29003.4]
  wire  _T_8881; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29004.4]
  wire  _T_8883; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29006.4]
  wire  _T_8884; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29007.4]
  wire  _T_8895; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29024.4]
  wire  _T_8896; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29025.4]
  wire  _T_8898; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29027.4]
  wire  _T_8900; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29029.4]
  wire [1:0] _T_8901; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29030.4]
  wire [1:0] _T_8902; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29031.4]
  wire  _T_8903; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29032.4]
  wire  _T_8904; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29034.4]
  wire  _T_8906; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29036.4]
  wire  _T_8908; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29038.4]
  wire  _T_8909; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29039.4]
  wire  _T_8910; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29044.4]
  wire  _T_8911; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29045.4]
  wire  _T_8912; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29046.4]
  wire  _T_8914; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29048.4]
  wire  _T_8915; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29049.4]
  wire  _T_8926; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29066.4]
  wire  _T_8927; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29067.4]
  wire  _T_8929; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29069.4]
  wire  _T_8931; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29071.4]
  wire [1:0] _T_8932; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29072.4]
  wire [1:0] _T_8933; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29073.4]
  wire  _T_8934; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29074.4]
  wire  _T_8935; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29076.4]
  wire  _T_8937; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29078.4]
  wire  _T_8939; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29080.4]
  wire  _T_8940; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29081.4]
  wire  _T_8941; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29086.4]
  wire  _T_8942; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29087.4]
  wire  _T_8943; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29088.4]
  wire  _T_8945; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29090.4]
  wire  _T_8946; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29091.4]
  wire  _T_8957; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29108.4]
  wire  _T_8958; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29109.4]
  wire  _T_8960; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29111.4]
  wire  _T_8962; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29113.4]
  wire [1:0] _T_8963; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29114.4]
  wire [1:0] _T_8964; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29115.4]
  wire  _T_8965; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29116.4]
  wire  _T_8966; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29118.4]
  wire  _T_8968; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29120.4]
  wire  _T_8970; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29122.4]
  wire  _T_8971; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29123.4]
  wire  _T_8972; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29128.4]
  wire  _T_8973; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29129.4]
  wire  _T_8974; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29130.4]
  wire  _T_8976; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29132.4]
  wire  _T_8977; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29133.4]
  wire  _T_8988; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29150.4]
  wire  _T_8989; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29151.4]
  wire  _T_8991; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29153.4]
  wire  _T_8993; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29155.4]
  wire [1:0] _T_8994; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29156.4]
  wire [1:0] _T_8995; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29157.4]
  wire  _T_8996; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29158.4]
  wire  _T_8997; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29160.4]
  wire  _T_8999; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29162.4]
  wire  _T_9001; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29164.4]
  wire  _T_9002; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29165.4]
  wire  _T_9003; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29170.4]
  wire  _T_9004; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29171.4]
  wire  _T_9005; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29172.4]
  wire  _T_9007; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29174.4]
  wire  _T_9008; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29175.4]
  wire  _T_9019; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29192.4]
  wire  _T_9020; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29193.4]
  wire  _T_9022; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29195.4]
  wire  _T_9024; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29197.4]
  wire [1:0] _T_9025; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29198.4]
  wire [1:0] _T_9026; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29199.4]
  wire  _T_9027; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29200.4]
  wire  _T_9028; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29202.4]
  wire  _T_9030; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29204.4]
  wire  _T_9032; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29206.4]
  wire  _T_9033; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29207.4]
  wire  _T_9034; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29212.4]
  wire  _T_9035; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29213.4]
  wire  _T_9036; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29214.4]
  wire  _T_9038; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29216.4]
  wire  _T_9039; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29217.4]
  wire  _T_9050; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29234.4]
  wire  _T_9051; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29235.4]
  wire  _T_9053; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29237.4]
  wire  _T_9055; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29239.4]
  wire [1:0] _T_9056; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29240.4]
  wire [1:0] _T_9057; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29241.4]
  wire  _T_9058; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29242.4]
  wire  _T_9059; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29244.4]
  wire  _T_9061; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29246.4]
  wire  _T_9063; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29248.4]
  wire  _T_9064; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29249.4]
  wire  _T_9065; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29254.4]
  wire  _T_9066; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29255.4]
  wire  _T_9067; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29256.4]
  wire  _T_9069; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29258.4]
  wire  _T_9070; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29259.4]
  wire  _T_9081; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29276.4]
  wire  _T_9082; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29277.4]
  wire  _T_9084; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29279.4]
  wire  _T_9086; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29281.4]
  wire [1:0] _T_9087; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29282.4]
  wire [1:0] _T_9088; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29283.4]
  wire  _T_9089; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29284.4]
  wire  _T_9090; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29286.4]
  wire  _T_9092; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29288.4]
  wire  _T_9094; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29290.4]
  wire  _T_9095; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29291.4]
  wire  _T_9096; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29296.4]
  wire  _T_9097; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29297.4]
  wire  _T_9098; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29298.4]
  wire  _T_9100; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29300.4]
  wire  _T_9101; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29301.4]
  wire  _T_9112; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29318.4]
  wire  _T_9113; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29319.4]
  wire  _T_9115; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29321.4]
  wire  _T_9117; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29323.4]
  wire [1:0] _T_9118; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29324.4]
  wire [1:0] _T_9119; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29325.4]
  wire  _T_9120; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29326.4]
  wire  _T_9121; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29328.4]
  wire  _T_9123; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29330.4]
  wire  _T_9125; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29332.4]
  wire  _T_9126; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29333.4]
  wire  _T_9127; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29338.4]
  wire  _T_9128; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29339.4]
  wire  _T_9129; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29340.4]
  wire  _T_9131; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29342.4]
  wire  _T_9132; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29343.4]
  wire  _T_9143; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29360.4]
  wire  _T_9144; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29361.4]
  wire  _T_9146; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29363.4]
  wire  _T_9148; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29365.4]
  wire [1:0] _T_9149; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29366.4]
  wire [1:0] _T_9150; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29367.4]
  wire  _T_9151; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29368.4]
  wire  _T_9152; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29370.4]
  wire  _T_9154; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29372.4]
  wire  _T_9156; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29374.4]
  wire  _T_9157; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29375.4]
  wire  _T_9158; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29380.4]
  wire  _T_9159; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29381.4]
  wire  _T_9160; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29382.4]
  wire  _T_9162; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29384.4]
  wire  _T_9163; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29385.4]
  wire  _T_9174; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29402.4]
  wire  _T_9175; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29403.4]
  wire  _T_9177; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29405.4]
  wire  _T_9179; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29407.4]
  wire [1:0] _T_9180; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29408.4]
  wire [1:0] _T_9181; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29409.4]
  wire  _T_9182; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29410.4]
  wire  _T_9183; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29412.4]
  wire  _T_9185; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29414.4]
  wire  _T_9187; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29416.4]
  wire  _T_9188; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29417.4]
  wire  _T_9189; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29422.4]
  wire  _T_9190; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29423.4]
  wire  _T_9191; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29424.4]
  wire  _T_9193; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29426.4]
  wire  _T_9194; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29427.4]
  wire  _T_9205; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29444.4]
  wire  _T_9206; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29445.4]
  wire  _T_9208; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29447.4]
  wire  _T_9210; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29449.4]
  wire [1:0] _T_9211; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29450.4]
  wire [1:0] _T_9212; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29451.4]
  wire  _T_9213; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29452.4]
  wire  _T_9214; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29454.4]
  wire  _T_9216; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29456.4]
  wire  _T_9218; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29458.4]
  wire  _T_9219; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29459.4]
  wire  _T_9220; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29464.4]
  wire  _T_9221; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29465.4]
  wire  _T_9222; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29466.4]
  wire  _T_9224; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29468.4]
  wire  _T_9225; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29469.4]
  wire  _T_9236; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29486.4]
  wire  _T_9237; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29487.4]
  wire  _T_9239; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29489.4]
  wire  _T_9241; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29491.4]
  wire [1:0] _T_9242; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29492.4]
  wire [1:0] _T_9243; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29493.4]
  wire  _T_9244; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29494.4]
  wire  _T_9245; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29496.4]
  wire  _T_9247; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29498.4]
  wire  _T_9249; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29500.4]
  wire  _T_9250; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29501.4]
  wire  _T_9251; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29506.4]
  wire  _T_9252; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29507.4]
  wire  _T_9253; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29508.4]
  wire  _T_9255; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29510.4]
  wire  _T_9256; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29511.4]
  wire  _T_9267; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29528.4]
  wire  _T_9268; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29529.4]
  wire  _T_9270; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29531.4]
  wire  _T_9272; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29533.4]
  wire [1:0] _T_9273; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29534.4]
  wire [1:0] _T_9274; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29535.4]
  wire  _T_9275; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29536.4]
  wire  _T_9276; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29538.4]
  wire  _T_9278; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29540.4]
  wire  _T_9280; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29542.4]
  wire  _T_9281; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29543.4]
  wire  _T_9282; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29548.4]
  wire  _T_9283; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29549.4]
  wire  _T_9284; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29550.4]
  wire  _T_9286; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29552.4]
  wire  _T_9287; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29553.4]
  wire  _T_9298; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29570.4]
  wire  _T_9299; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29571.4]
  wire  _T_9301; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29573.4]
  wire  _T_9303; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29575.4]
  wire [1:0] _T_9304; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29576.4]
  wire [1:0] _T_9305; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29577.4]
  wire  _T_9306; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29578.4]
  wire  _T_9307; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29580.4]
  wire  _T_9309; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29582.4]
  wire  _T_9311; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29584.4]
  wire  _T_9312; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29585.4]
  wire  _T_9313; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29590.4]
  wire  _T_9314; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29591.4]
  wire  _T_9315; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29592.4]
  wire  _T_9317; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29594.4]
  wire  _T_9318; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29595.4]
  wire  _T_9329; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29612.4]
  wire  _T_9330; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29613.4]
  wire  _T_9332; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29615.4]
  wire  _T_9334; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29617.4]
  wire [1:0] _T_9335; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29618.4]
  wire [1:0] _T_9336; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29619.4]
  wire  _T_9337; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29620.4]
  wire  _T_9338; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29622.4]
  wire  _T_9340; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29624.4]
  wire  _T_9342; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29626.4]
  wire  _T_9343; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29627.4]
  wire  _T_9344; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29632.4]
  wire  _T_9345; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29633.4]
  wire  _T_9346; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29634.4]
  wire  _T_9348; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29636.4]
  wire  _T_9349; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29637.4]
  wire  _T_9360; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29654.4]
  wire  _T_9361; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29655.4]
  wire  _T_9363; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29657.4]
  wire  _T_9365; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29659.4]
  wire [1:0] _T_9366; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29660.4]
  wire [1:0] _T_9367; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29661.4]
  wire  _T_9368; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29662.4]
  wire  _T_9369; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29664.4]
  wire  _T_9371; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29666.4]
  wire  _T_9373; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29668.4]
  wire  _T_9374; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29669.4]
  wire  _T_9375; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29674.4]
  wire  _T_9376; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29675.4]
  wire  _T_9377; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29676.4]
  wire  _T_9379; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29678.4]
  wire  _T_9380; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29679.4]
  wire  _T_9391; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29696.4]
  wire  _T_9392; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29697.4]
  wire  _T_9394; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29699.4]
  wire  _T_9396; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29701.4]
  wire [1:0] _T_9397; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29702.4]
  wire [1:0] _T_9398; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29703.4]
  wire  _T_9399; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29704.4]
  wire  _T_9400; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29706.4]
  wire  _T_9402; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29708.4]
  wire  _T_9404; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29710.4]
  wire  _T_9405; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29711.4]
  wire  _T_9406; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29716.4]
  wire  _T_9407; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29717.4]
  wire  _T_9408; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29718.4]
  wire  _T_9410; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29720.4]
  wire  _T_9411; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29721.4]
  wire  _T_9422; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29738.4]
  wire  _T_9423; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29739.4]
  wire  _T_9425; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29741.4]
  wire  _T_9427; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29743.4]
  wire [1:0] _T_9428; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29744.4]
  wire [1:0] _T_9429; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29745.4]
  wire  _T_9430; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29746.4]
  wire  _T_9431; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29748.4]
  wire  _T_9433; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29750.4]
  wire  _T_9435; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29752.4]
  wire  _T_9436; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29753.4]
  wire  _T_9437; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29758.4]
  wire  _T_9438; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29759.4]
  wire  _T_9439; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29760.4]
  wire  _T_9441; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29762.4]
  wire  _T_9442; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29763.4]
  wire  _T_9453; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29780.4]
  wire  _T_9454; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29781.4]
  wire  _T_9456; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29783.4]
  wire  _T_9458; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29785.4]
  wire [1:0] _T_9459; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29786.4]
  wire [1:0] _T_9460; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29787.4]
  wire  _T_9461; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29788.4]
  wire  _T_9462; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29790.4]
  wire  _T_9464; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29792.4]
  wire  _T_9466; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29794.4]
  wire  _T_9467; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29795.4]
  wire  _T_9468; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29800.4]
  wire  _T_9469; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29801.4]
  wire  _T_9470; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29802.4]
  wire  _T_9472; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29804.4]
  wire  _T_9473; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29805.4]
  wire  _T_9484; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29822.4]
  wire  _T_9485; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29823.4]
  wire  _T_9487; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29825.4]
  wire  _T_9489; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29827.4]
  wire [1:0] _T_9490; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29828.4]
  wire [1:0] _T_9491; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29829.4]
  wire  _T_9492; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29830.4]
  wire  _T_9493; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29832.4]
  wire  _T_9495; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29834.4]
  wire  _T_9497; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29836.4]
  wire  _T_9498; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29837.4]
  wire  _T_9499; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29842.4]
  wire  _T_9500; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29843.4]
  wire  _T_9501; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29844.4]
  wire  _T_9503; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29846.4]
  wire  _T_9504; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29847.4]
  wire  _T_9515; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29864.4]
  wire  _T_9516; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29865.4]
  wire  _T_9518; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29867.4]
  wire  _T_9520; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29869.4]
  wire [1:0] _T_9521; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29870.4]
  wire [1:0] _T_9522; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29871.4]
  wire  _T_9523; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29872.4]
  wire  _T_9524; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29874.4]
  wire  _T_9526; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29876.4]
  wire  _T_9528; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29878.4]
  wire  _T_9529; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29879.4]
  wire  _T_9530; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29884.4]
  wire  _T_9531; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29885.4]
  wire  _T_9532; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29886.4]
  wire  _T_9534; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29888.4]
  wire  _T_9535; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29889.4]
  wire  _T_9546; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29906.4]
  wire  _T_9547; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29907.4]
  wire  _T_9549; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29909.4]
  wire  _T_9551; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29911.4]
  wire [1:0] _T_9552; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29912.4]
  wire [1:0] _T_9553; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29913.4]
  wire  _T_9554; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29914.4]
  wire  _T_9555; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29916.4]
  wire  _T_9557; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29918.4]
  wire  _T_9559; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29920.4]
  wire  _T_9560; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29921.4]
  wire  _T_9561; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29926.4]
  wire  _T_9562; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29927.4]
  wire  _T_9563; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29928.4]
  wire  _T_9565; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29930.4]
  wire  _T_9566; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29931.4]
  wire  _T_9577; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29948.4]
  wire  _T_9578; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29949.4]
  wire  _T_9580; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29951.4]
  wire  _T_9582; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29953.4]
  wire [1:0] _T_9583; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29954.4]
  wire [1:0] _T_9584; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29955.4]
  wire  _T_9585; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29956.4]
  wire  _T_9586; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29958.4]
  wire  _T_9588; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29960.4]
  wire  _T_9590; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29962.4]
  wire  _T_9591; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29963.4]
  wire  _T_9592; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29968.4]
  wire  _T_9593; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29969.4]
  wire  _T_9594; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29970.4]
  wire  _T_9596; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29972.4]
  wire  _T_9597; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29973.4]
  wire  _T_9608; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29990.4]
  wire  _T_9609; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29991.4]
  wire  _T_9611; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29993.4]
  wire  _T_9613; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29995.4]
  wire [1:0] _T_9614; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29996.4]
  wire [1:0] _T_9615; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29997.4]
  wire  _T_9616; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29998.4]
  wire  _T_9617; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30000.4]
  wire  _T_9619; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30002.4]
  wire  _T_9621; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30004.4]
  wire  _T_9622; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30005.4]
  wire  _T_9623; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30010.4]
  wire  _T_9624; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30011.4]
  wire  _T_9625; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30012.4]
  wire  _T_9627; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30014.4]
  wire  _T_9628; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30015.4]
  wire  _T_9639; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30032.4]
  wire  _T_9640; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30033.4]
  wire  _T_9642; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30035.4]
  wire  _T_9644; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30037.4]
  wire [1:0] _T_9645; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30038.4]
  wire [1:0] _T_9646; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30039.4]
  wire  _T_9647; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30040.4]
  wire  _T_9648; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30042.4]
  wire  _T_9650; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30044.4]
  wire  _T_9652; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30046.4]
  wire  _T_9653; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30047.4]
  wire  _T_9654; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30052.4]
  wire  _T_9655; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30053.4]
  wire  _T_9656; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30054.4]
  wire  _T_9658; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30056.4]
  wire  _T_9659; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30057.4]
  wire  _T_9670; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30074.4]
  wire  _T_9671; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30075.4]
  wire  _T_9673; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30077.4]
  wire  _T_9675; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30079.4]
  wire [1:0] _T_9676; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30080.4]
  wire [1:0] _T_9677; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30081.4]
  wire  _T_9678; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30082.4]
  wire  _T_9679; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30084.4]
  wire  _T_9681; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30086.4]
  wire  _T_9683; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30088.4]
  wire  _T_9684; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30089.4]
  wire  _T_9685; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30094.4]
  wire  _T_9686; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30095.4]
  wire  _T_9687; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30096.4]
  wire  _T_9689; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30098.4]
  wire  _T_9690; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30099.4]
  wire  _T_9701; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30116.4]
  wire  _T_9702; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30117.4]
  wire  _T_9704; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30119.4]
  wire  _T_9706; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30121.4]
  wire [1:0] _T_9707; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30122.4]
  wire [1:0] _T_9708; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30123.4]
  wire  _T_9709; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30124.4]
  wire  _T_9710; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30126.4]
  wire  _T_9712; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30128.4]
  wire  _T_9714; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30130.4]
  wire  _T_9715; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30131.4]
  wire  _T_9716; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30136.4]
  wire  _T_9717; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30137.4]
  wire  _T_9718; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30138.4]
  wire  _T_9720; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30140.4]
  wire  _T_9721; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30141.4]
  wire  _T_9732; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30158.4]
  wire  _T_9733; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30159.4]
  wire  _T_9735; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30161.4]
  wire  _T_9737; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30163.4]
  wire [1:0] _T_9738; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30164.4]
  wire [1:0] _T_9739; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30165.4]
  wire  _T_9740; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30166.4]
  wire  _T_9741; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30168.4]
  wire  _T_9743; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30170.4]
  wire  _T_9745; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30172.4]
  wire  _T_9746; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30173.4]
  wire  _T_9747; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30178.4]
  wire  _T_9748; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30179.4]
  wire  _T_9749; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30180.4]
  wire  _T_9751; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30182.4]
  wire  _T_9752; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30183.4]
  wire  _T_9763; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30200.4]
  wire  _T_9764; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30201.4]
  wire  _T_9766; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30203.4]
  wire  _T_9768; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30205.4]
  wire [1:0] _T_9769; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30206.4]
  wire [1:0] _T_9770; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30207.4]
  wire  _T_9771; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30208.4]
  wire  _T_9772; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30210.4]
  wire  _T_9774; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30212.4]
  wire  _T_9776; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30214.4]
  wire  _T_9777; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30215.4]
  wire  _T_9778; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30220.4]
  wire  _T_9779; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30221.4]
  wire  _T_9780; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30222.4]
  wire  _T_9782; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30224.4]
  wire  _T_9783; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30225.4]
  wire  _T_9794; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30242.4]
  wire  _T_9795; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30243.4]
  wire  _T_9797; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30245.4]
  wire  _T_9799; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30247.4]
  wire [1:0] _T_9800; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30248.4]
  wire [1:0] _T_9801; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30249.4]
  wire  _T_9802; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30250.4]
  wire  _T_9803; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30252.4]
  wire  _T_9805; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30254.4]
  wire  _T_9807; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30256.4]
  wire  _T_9808; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30257.4]
  wire  _T_9809; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30262.4]
  wire  _T_9810; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30263.4]
  wire  _T_9811; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30264.4]
  wire  _T_9813; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30266.4]
  wire  _T_9814; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30267.4]
  wire  _T_9825; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30284.4]
  wire  _T_9826; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30285.4]
  wire  _T_9828; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30287.4]
  wire  _T_9830; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30289.4]
  wire [1:0] _T_9831; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30290.4]
  wire [1:0] _T_9832; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30291.4]
  wire  _T_9833; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30292.4]
  wire  _T_9834; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30294.4]
  wire  _T_9836; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30296.4]
  wire  _T_9838; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30298.4]
  wire  _T_9839; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30299.4]
  wire  _T_9840; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30304.4]
  wire  _T_9841; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30305.4]
  wire  _T_9842; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30306.4]
  wire  _T_9844; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30308.4]
  wire  _T_9845; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30309.4]
  wire  _T_9856; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30326.4]
  wire  _T_9857; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30327.4]
  wire  _T_9859; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30329.4]
  wire  _T_9861; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30331.4]
  wire [1:0] _T_9862; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30332.4]
  wire [1:0] _T_9863; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30333.4]
  wire  _T_9864; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30334.4]
  wire  _T_9865; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30336.4]
  wire  _T_9867; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30338.4]
  wire  _T_9869; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30340.4]
  wire  _T_9870; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30341.4]
  wire  _T_9871; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30346.4]
  wire  _T_9872; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30347.4]
  wire  _T_9873; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30348.4]
  wire  _T_9875; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30350.4]
  wire  _T_9876; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30351.4]
  wire  _T_9887; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30368.4]
  wire  _T_9888; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30369.4]
  wire  _T_9890; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30371.4]
  wire  _T_9892; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30373.4]
  wire [1:0] _T_9893; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30374.4]
  wire [1:0] _T_9894; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30375.4]
  wire  _T_9895; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30376.4]
  wire  _T_9896; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30378.4]
  wire  _T_9898; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30380.4]
  wire  _T_9900; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30382.4]
  wire  _T_9901; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30383.4]
  wire  _T_9902; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30388.4]
  wire  _T_9903; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30389.4]
  wire  _T_9904; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30390.4]
  wire  _T_9906; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30392.4]
  wire  _T_9907; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30393.4]
  wire  _T_9918; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30410.4]
  wire  _T_9919; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30411.4]
  wire  _T_9921; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30413.4]
  wire  _T_9923; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30415.4]
  wire [1:0] _T_9924; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30416.4]
  wire [1:0] _T_9925; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30417.4]
  wire  _T_9926; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30418.4]
  wire  _T_9927; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30420.4]
  wire  _T_9929; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30422.4]
  wire  _T_9931; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30424.4]
  wire  _T_9932; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30425.4]
  wire  _T_9933; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30430.4]
  wire  _T_9934; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30431.4]
  wire  _T_9935; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30432.4]
  wire  _T_9937; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30434.4]
  wire  _T_9938; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30435.4]
  wire  _T_9949; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30452.4]
  wire  _T_9950; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30453.4]
  wire  _T_9952; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30455.4]
  wire  _T_9954; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30457.4]
  wire [1:0] _T_9955; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30458.4]
  wire [1:0] _T_9956; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30459.4]
  wire  _T_9957; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30460.4]
  wire  _T_9958; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30462.4]
  wire  _T_9960; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30464.4]
  wire  _T_9962; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30466.4]
  wire  _T_9963; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30467.4]
  wire  _T_9964; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30472.4]
  wire  _T_9965; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30473.4]
  wire  _T_9966; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30474.4]
  wire  _T_9968; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30476.4]
  wire  _T_9969; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30477.4]
  wire  _T_9980; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30494.4]
  wire  _T_9981; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30495.4]
  wire  _T_9983; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30497.4]
  wire  _T_9985; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30499.4]
  wire [1:0] _T_9986; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30500.4]
  wire [1:0] _T_9987; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30501.4]
  wire  _T_9988; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30502.4]
  wire  _T_9989; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30504.4]
  wire  _T_9991; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30506.4]
  wire  _T_9993; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30508.4]
  wire  _T_9994; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30509.4]
  wire  _T_9995; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30514.4]
  wire  _T_9996; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30515.4]
  wire  _T_9997; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30516.4]
  wire  _T_9999; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30518.4]
  wire  _T_10000; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30519.4]
  wire  _T_10011; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30536.4]
  wire  _T_10012; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30537.4]
  wire  _T_10014; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30539.4]
  wire  _T_10016; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30541.4]
  wire [1:0] _T_10017; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30542.4]
  wire [1:0] _T_10018; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30543.4]
  wire  _T_10019; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30544.4]
  wire  _T_10020; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30546.4]
  wire  _T_10022; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30548.4]
  wire  _T_10024; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30550.4]
  wire  _T_10025; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30551.4]
  wire  _T_10026; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30556.4]
  wire  _T_10027; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30557.4]
  wire  _T_10028; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30558.4]
  wire  _T_10030; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30560.4]
  wire  _T_10031; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30561.4]
  wire  _T_10042; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30578.4]
  wire  _T_10043; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30579.4]
  wire  _T_10045; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30581.4]
  wire  _T_10047; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30583.4]
  wire [1:0] _T_10048; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30584.4]
  wire [1:0] _T_10049; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30585.4]
  wire  _T_10050; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30586.4]
  wire  _T_10051; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30588.4]
  wire  _T_10053; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30590.4]
  wire  _T_10055; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30592.4]
  wire  _T_10056; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30593.4]
  wire  _T_10057; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30598.4]
  wire  _T_10058; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30599.4]
  wire  _T_10059; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30600.4]
  wire  _T_10061; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30602.4]
  wire  _T_10062; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30603.4]
  wire  _T_10073; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30620.4]
  wire  _T_10074; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30621.4]
  wire  _T_10076; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30623.4]
  wire  _T_10078; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30625.4]
  wire [1:0] _T_10079; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30626.4]
  wire [1:0] _T_10080; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30627.4]
  wire  _T_10081; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30628.4]
  wire  _T_10082; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30630.4]
  wire  _T_10084; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30632.4]
  wire  _T_10086; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30634.4]
  wire  _T_10087; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30635.4]
  wire  _T_10088; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30640.4]
  wire  _T_10089; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30641.4]
  wire  _T_10090; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30642.4]
  wire  _T_10092; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30644.4]
  wire  _T_10093; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30645.4]
  wire  _T_10104; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30662.4]
  wire  _T_10105; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30663.4]
  wire  _T_10107; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30665.4]
  wire  _T_10109; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30667.4]
  wire [1:0] _T_10110; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30668.4]
  wire [1:0] _T_10111; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30669.4]
  wire  _T_10112; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30670.4]
  wire  _T_10113; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30672.4]
  wire  _T_10115; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30674.4]
  wire  _T_10117; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30676.4]
  wire  _T_10118; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30677.4]
  wire  _T_10119; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30682.4]
  wire  _T_10120; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30683.4]
  wire  _T_10121; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30684.4]
  wire  _T_10123; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30686.4]
  wire  _T_10124; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30687.4]
  wire  _T_10135; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30704.4]
  wire  _T_10136; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30705.4]
  wire  _T_10138; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30707.4]
  wire  _T_10140; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30709.4]
  wire [1:0] _T_10141; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30710.4]
  wire [1:0] _T_10142; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30711.4]
  wire  _T_10143; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30712.4]
  wire  _T_10144; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30714.4]
  wire  _T_10146; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30716.4]
  wire  _T_10148; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30718.4]
  wire  _T_10149; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30719.4]
  wire  _T_10150; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30724.4]
  wire  _T_10151; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30725.4]
  wire  _T_10152; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30726.4]
  wire  _T_10154; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30728.4]
  wire  _T_10155; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30729.4]
  wire  _T_10166; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30746.4]
  wire  _T_10167; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30747.4]
  wire  _T_10169; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30749.4]
  wire  _T_10171; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30751.4]
  wire [1:0] _T_10172; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30752.4]
  wire [1:0] _T_10173; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30753.4]
  wire  _T_10174; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30754.4]
  wire  _T_10175; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30756.4]
  wire  _T_10177; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30758.4]
  wire  _T_10179; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30760.4]
  wire  _T_10180; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30761.4]
  wire  _T_10181; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30766.4]
  wire  _T_10182; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30767.4]
  wire  _T_10183; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30768.4]
  wire  _T_10185; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30770.4]
  wire  _T_10186; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30771.4]
  wire  _T_10197; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30788.4]
  wire  _T_10198; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30789.4]
  wire  _T_10200; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30791.4]
  wire  _T_10202; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30793.4]
  wire [1:0] _T_10203; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30794.4]
  wire [1:0] _T_10204; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30795.4]
  wire  _T_10205; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30796.4]
  wire  _T_10206; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30798.4]
  wire  _T_10208; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30800.4]
  wire  _T_10210; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30802.4]
  wire  _T_10211; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30803.4]
  wire  _T_10212; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30808.4]
  wire  _T_10213; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30809.4]
  wire  _T_10214; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30810.4]
  wire  _T_10216; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30812.4]
  wire  _T_10217; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30813.4]
  wire  _T_10228; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30830.4]
  wire  _T_10229; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30831.4]
  wire  _T_10231; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30833.4]
  wire  _T_10233; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30835.4]
  wire [1:0] _T_10234; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30836.4]
  wire [1:0] _T_10235; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30837.4]
  wire  _T_10236; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30838.4]
  wire  _T_10237; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30840.4]
  wire  _T_10239; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30842.4]
  wire  _T_10241; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30844.4]
  wire  _T_10242; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30845.4]
  wire  _T_10243; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30850.4]
  wire  _T_10244; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30851.4]
  wire  _T_10245; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30852.4]
  wire  _T_10247; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30854.4]
  wire  _T_10248; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30855.4]
  wire  _T_10259; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30872.4]
  wire  _T_10260; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30873.4]
  wire  _T_10262; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30875.4]
  wire  _T_10264; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30877.4]
  wire [1:0] _T_10265; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30878.4]
  wire [1:0] _T_10266; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30879.4]
  wire  _T_10267; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30880.4]
  wire  _T_10268; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30882.4]
  wire  _T_10270; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30884.4]
  wire  _T_10272; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30886.4]
  wire  _T_10273; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30887.4]
  wire  _T_10274; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30892.4]
  wire  _T_10275; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30893.4]
  wire  _T_10276; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30894.4]
  wire  _T_10278; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30896.4]
  wire  _T_10279; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30897.4]
  wire  _T_10290; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30914.4]
  wire  _T_10291; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30915.4]
  wire  _T_10293; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30917.4]
  wire  _T_10295; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30919.4]
  wire [1:0] _T_10296; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30920.4]
  wire [1:0] _T_10297; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30921.4]
  wire  _T_10298; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30922.4]
  wire  _T_10299; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30924.4]
  wire  _T_10301; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30926.4]
  wire  _T_10303; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30928.4]
  wire  _T_10304; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30929.4]
  wire  _T_10305; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30934.4]
  wire  _T_10306; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30935.4]
  wire  _T_10307; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30936.4]
  wire  _T_10309; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30938.4]
  wire  _T_10310; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30939.4]
  wire  _T_10321; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30956.4]
  wire  _T_10322; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30957.4]
  wire  _T_10324; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30959.4]
  wire  _T_10326; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30961.4]
  wire [1:0] _T_10327; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30962.4]
  wire [1:0] _T_10328; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30963.4]
  wire  _T_10329; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30964.4]
  wire  _T_10330; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30966.4]
  wire  _T_10332; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30968.4]
  wire  _T_10334; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30970.4]
  wire  _T_10335; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30971.4]
  wire  _T_10336; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30976.4]
  wire  _T_10337; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30977.4]
  wire  _T_10338; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30978.4]
  wire  _T_10340; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30980.4]
  wire  _T_10341; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30981.4]
  wire  _T_10352; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30998.4]
  wire  _T_10353; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30999.4]
  wire  _T_10355; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31001.4]
  wire  _T_10357; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31003.4]
  wire [1:0] _T_10358; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31004.4]
  wire [1:0] _T_10359; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31005.4]
  wire  _T_10360; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31006.4]
  wire  _T_10361; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31008.4]
  wire  _T_10363; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31010.4]
  wire  _T_10365; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31012.4]
  wire  _T_10366; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31013.4]
  wire  _T_10367; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31018.4]
  wire  _T_10368; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31019.4]
  wire  _T_10369; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31020.4]
  wire  _T_10371; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31022.4]
  wire  _T_10372; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31023.4]
  wire  _T_10383; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31040.4]
  wire  _T_10384; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31041.4]
  wire  _T_10386; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31043.4]
  wire  _T_10388; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31045.4]
  wire [1:0] _T_10389; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31046.4]
  wire [1:0] _T_10390; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31047.4]
  wire  _T_10391; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31048.4]
  wire  _T_10392; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31050.4]
  wire  _T_10394; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31052.4]
  wire  _T_10396; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31054.4]
  wire  _T_10397; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31055.4]
  wire  _T_10398; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31060.4]
  wire  _T_10399; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31061.4]
  wire  _T_10400; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31062.4]
  wire  _T_10402; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31064.4]
  wire  _T_10403; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31065.4]
  wire  _T_10414; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31082.4]
  wire  _T_10415; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31083.4]
  wire  _T_10417; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31085.4]
  wire  _T_10419; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31087.4]
  wire [1:0] _T_10420; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31088.4]
  wire [1:0] _T_10421; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31089.4]
  wire  _T_10422; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31090.4]
  wire  _T_10423; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31092.4]
  wire  _T_10425; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31094.4]
  wire  _T_10427; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31096.4]
  wire  _T_10428; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31097.4]
  wire  _T_10429; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31102.4]
  wire  _T_10430; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31103.4]
  wire  _T_10431; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31104.4]
  wire  _T_10433; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31106.4]
  wire  _T_10434; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31107.4]
  wire  _T_10445; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31124.4]
  wire  _T_10446; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31125.4]
  wire  _T_10448; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31127.4]
  wire  _T_10450; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31129.4]
  wire [1:0] _T_10451; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31130.4]
  wire [1:0] _T_10452; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31131.4]
  wire  _T_10453; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31132.4]
  wire  _T_10454; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31134.4]
  wire  _T_10456; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31136.4]
  wire  _T_10458; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31138.4]
  wire  _T_10459; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31139.4]
  wire  _T_10460; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31144.4]
  wire  _T_10461; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31145.4]
  wire  _T_10462; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31146.4]
  wire  _T_10464; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31148.4]
  wire  _T_10465; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31149.4]
  wire  _T_10476; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31166.4]
  wire  _T_10477; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31167.4]
  wire  _T_10479; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31169.4]
  wire  _T_10481; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31171.4]
  wire [1:0] _T_10482; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31172.4]
  wire [1:0] _T_10483; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31173.4]
  wire  _T_10484; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31174.4]
  wire  _T_10485; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31176.4]
  wire  _T_10487; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31178.4]
  wire  _T_10489; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31180.4]
  wire  _T_10490; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31181.4]
  wire  _T_10491; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31186.4]
  wire  _T_10492; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31187.4]
  wire  _T_10493; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31188.4]
  wire  _T_10495; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31190.4]
  wire  _T_10496; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31191.4]
  wire  _T_10507; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31208.4]
  wire  _T_10508; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31209.4]
  wire  _T_10510; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31211.4]
  wire  _T_10512; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31213.4]
  wire [1:0] _T_10513; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31214.4]
  wire [1:0] _T_10514; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31215.4]
  wire  _T_10515; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31216.4]
  wire  _T_10516; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31218.4]
  wire  _T_10518; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31220.4]
  wire  _T_10520; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31222.4]
  wire  _T_10521; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31223.4]
  wire  _T_10522; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31228.4]
  wire  _T_10523; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31229.4]
  wire  _T_10524; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31230.4]
  wire  _T_10526; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31232.4]
  wire  _T_10527; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31233.4]
  wire  _T_10538; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31250.4]
  wire  _T_10539; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31251.4]
  wire  _T_10541; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31253.4]
  wire  _T_10543; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31255.4]
  wire [1:0] _T_10544; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31256.4]
  wire [1:0] _T_10545; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31257.4]
  wire  _T_10546; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31258.4]
  wire  _T_10547; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31260.4]
  wire  _T_10549; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31262.4]
  wire  _T_10551; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31264.4]
  wire  _T_10552; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31265.4]
  wire  _T_10553; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31270.4]
  wire  _T_10554; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31271.4]
  wire  _T_10555; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31272.4]
  wire  _T_10557; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31274.4]
  wire  _T_10558; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31275.4]
  wire  _T_10569; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31292.4]
  wire  _T_10570; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31293.4]
  wire  _T_10572; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31295.4]
  wire  _T_10574; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31297.4]
  wire [1:0] _T_10575; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31298.4]
  wire [1:0] _T_10576; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31299.4]
  wire  _T_10577; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31300.4]
  wire  _T_10578; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31302.4]
  wire  _T_10580; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31304.4]
  wire  _T_10582; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31306.4]
  wire  _T_10583; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31307.4]
  wire  _T_10584; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31312.4]
  wire  _T_10585; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31313.4]
  wire  _T_10586; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31314.4]
  wire  _T_10588; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31316.4]
  wire  _T_10589; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31317.4]
  wire  _T_10600; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31334.4]
  wire  _T_10601; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31335.4]
  wire  _T_10603; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31337.4]
  wire  _T_10605; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31339.4]
  wire [1:0] _T_10606; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31340.4]
  wire [1:0] _T_10607; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31341.4]
  wire  _T_10608; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31342.4]
  wire  _T_10609; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31344.4]
  wire  _T_10611; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31346.4]
  wire  _T_10613; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31348.4]
  wire  _T_10614; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31349.4]
  wire  _T_10615; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31354.4]
  wire  _T_10616; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31355.4]
  wire  _T_10617; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31356.4]
  wire  _T_10619; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31358.4]
  wire  _T_10620; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31359.4]
  wire  _T_10631; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31376.4]
  wire  _T_10632; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31377.4]
  wire  _T_10634; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31379.4]
  wire  _T_10636; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31381.4]
  wire [1:0] _T_10637; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31382.4]
  wire [1:0] _T_10638; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31383.4]
  wire  _T_10639; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31384.4]
  wire  _T_10640; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31386.4]
  wire  _T_10642; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31388.4]
  wire  _T_10644; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31390.4]
  wire  _T_10645; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31391.4]
  wire  _T_10646; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31396.4]
  wire  _T_10647; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31397.4]
  wire  _T_10648; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31398.4]
  wire  _T_10650; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31400.4]
  wire  _T_10651; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31401.4]
  wire  _T_10662; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31418.4]
  wire  _T_10663; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31419.4]
  wire  _T_10665; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31421.4]
  wire  _T_10667; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31423.4]
  wire [1:0] _T_10668; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31424.4]
  wire [1:0] _T_10669; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31425.4]
  wire  _T_10670; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31426.4]
  wire  _T_10671; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31428.4]
  wire  _T_10673; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31430.4]
  wire  _T_10675; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31432.4]
  wire  _T_10676; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31433.4]
  wire  _T_10677; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31438.4]
  wire  _T_10678; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31439.4]
  wire  _T_10679; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31440.4]
  wire  _T_10681; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31442.4]
  wire  _T_10682; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31443.4]
  wire  _T_10693; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31460.4]
  wire  _T_10694; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31461.4]
  wire  _T_10696; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31463.4]
  wire  _T_10698; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31465.4]
  wire [1:0] _T_10699; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31466.4]
  wire [1:0] _T_10700; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31467.4]
  wire  _T_10701; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31468.4]
  wire  _T_10702; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31470.4]
  wire  _T_10704; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31472.4]
  wire  _T_10706; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31474.4]
  wire  _T_10707; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31475.4]
  wire  _T_10708; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31480.4]
  wire  _T_10709; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31481.4]
  wire  _T_10710; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31482.4]
  wire  _T_10712; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31484.4]
  wire  _T_10713; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31485.4]
  wire  _T_10724; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31502.4]
  wire  _T_10725; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31503.4]
  wire  _T_10727; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31505.4]
  wire  _T_10729; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31507.4]
  wire [1:0] _T_10730; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31508.4]
  wire [1:0] _T_10731; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31509.4]
  wire  _T_10732; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31510.4]
  wire  _T_10733; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31512.4]
  wire  _T_10735; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31514.4]
  wire  _T_10737; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31516.4]
  wire  _T_10738; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31517.4]
  wire  _T_10739; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31522.4]
  wire  _T_10740; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31523.4]
  wire  _T_10741; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31524.4]
  wire  _T_10743; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31526.4]
  wire  _T_10744; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31527.4]
  wire  _T_10755; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31544.4]
  wire  _T_10756; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31545.4]
  wire  _T_10758; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31547.4]
  wire  _T_10760; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31549.4]
  wire [1:0] _T_10761; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31550.4]
  wire [1:0] _T_10762; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31551.4]
  wire  _T_10763; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31552.4]
  wire  _T_10764; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31554.4]
  wire  _T_10766; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31556.4]
  wire  _T_10768; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31558.4]
  wire  _T_10769; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31559.4]
  wire  _T_10770; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31564.4]
  wire  _T_10771; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31565.4]
  wire  _T_10772; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31566.4]
  wire  _T_10774; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31568.4]
  wire  _T_10775; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31569.4]
  wire  _T_10786; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31586.4]
  wire  _T_10787; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31587.4]
  wire  _T_10789; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31589.4]
  wire  _T_10791; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31591.4]
  wire [1:0] _T_10792; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31592.4]
  wire [1:0] _T_10793; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31593.4]
  wire  _T_10794; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31594.4]
  wire  _T_10795; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31596.4]
  wire  _T_10797; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31598.4]
  wire  _T_10799; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31600.4]
  wire  _T_10800; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31601.4]
  wire  _T_10801; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31606.4]
  wire  _T_10802; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31607.4]
  wire  _T_10803; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31608.4]
  wire  _T_10805; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31610.4]
  wire  _T_10806; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31611.4]
  wire  _T_10817; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31628.4]
  wire  _T_10818; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31629.4]
  wire  _T_10820; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31631.4]
  wire  _T_10822; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31633.4]
  wire [1:0] _T_10823; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31634.4]
  wire [1:0] _T_10824; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31635.4]
  wire  _T_10825; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31636.4]
  wire  _T_10826; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31638.4]
  wire  _T_10828; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31640.4]
  wire  _T_10830; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31642.4]
  wire  _T_10831; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31643.4]
  wire  _T_10832; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31648.4]
  wire  _T_10833; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31649.4]
  wire  _T_10834; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31650.4]
  wire  _T_10836; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31652.4]
  wire  _T_10837; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31653.4]
  wire  _T_10848; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31670.4]
  wire  _T_10849; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31671.4]
  wire  _T_10851; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31673.4]
  wire  _T_10853; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31675.4]
  wire [1:0] _T_10854; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31676.4]
  wire [1:0] _T_10855; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31677.4]
  wire  _T_10856; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31678.4]
  wire  _T_10857; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31680.4]
  wire  _T_10859; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31682.4]
  wire  _T_10861; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31684.4]
  wire  _T_10862; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31685.4]
  wire  _T_10863; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31690.4]
  wire  _T_10864; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31691.4]
  wire  _T_10865; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31692.4]
  wire  _T_10867; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31694.4]
  wire  _T_10868; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31695.4]
  Queue_43 Queue ( // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20285.4]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_strb(Queue_io_enq_bits_strb),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_strb(Queue_io_deq_bits_strb),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_97 Queue_1 ( // @[Decoupled.scala 293:21:boom.system.TestHarness.MegaBoomConfig.fir@20300.4]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_wen(Queue_1_io_enq_bits_wen),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_1_io_deq_bits_qos),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_wen(Queue_1_io_deq_bits_wen)
  );
  assign _T_2295 = auto_in_a_bits_opcode[2]; // @[Edges.scala 92:37:boom.system.TestHarness.MegaBoomConfig.fir@20232.4]
  assign _T_2296 = _T_2295 == 1'h0; // @[Edges.scala 92:28:boom.system.TestHarness.MegaBoomConfig.fir@20233.4]
  assign _GEN_259 = 8'h1 == auto_in_a_bits_source ? _T_2969 : _T_2938; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_260 = 8'h2 == auto_in_a_bits_source ? _T_3000 : _GEN_259; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_261 = 8'h3 == auto_in_a_bits_source ? _T_3031 : _GEN_260; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_262 = 8'h4 == auto_in_a_bits_source ? _T_3062 : _GEN_261; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_263 = 8'h5 == auto_in_a_bits_source ? _T_3093 : _GEN_262; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_264 = 8'h6 == auto_in_a_bits_source ? _T_3124 : _GEN_263; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_265 = 8'h7 == auto_in_a_bits_source ? _T_3155 : _GEN_264; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_266 = 8'h8 == auto_in_a_bits_source ? _T_3186 : _GEN_265; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_267 = 8'h9 == auto_in_a_bits_source ? _T_3217 : _GEN_266; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_268 = 8'ha == auto_in_a_bits_source ? _T_3248 : _GEN_267; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_269 = 8'hb == auto_in_a_bits_source ? _T_3279 : _GEN_268; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_270 = 8'hc == auto_in_a_bits_source ? _T_3310 : _GEN_269; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_271 = 8'hd == auto_in_a_bits_source ? _T_3341 : _GEN_270; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_272 = 8'he == auto_in_a_bits_source ? _T_3372 : _GEN_271; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_273 = 8'hf == auto_in_a_bits_source ? _T_3403 : _GEN_272; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_274 = 8'h10 == auto_in_a_bits_source ? _T_3434 : _GEN_273; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_275 = 8'h11 == auto_in_a_bits_source ? _T_3465 : _GEN_274; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_276 = 8'h12 == auto_in_a_bits_source ? _T_3496 : _GEN_275; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_277 = 8'h13 == auto_in_a_bits_source ? _T_3527 : _GEN_276; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_278 = 8'h14 == auto_in_a_bits_source ? _T_3558 : _GEN_277; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_279 = 8'h15 == auto_in_a_bits_source ? _T_3589 : _GEN_278; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_280 = 8'h16 == auto_in_a_bits_source ? _T_3620 : _GEN_279; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_281 = 8'h17 == auto_in_a_bits_source ? _T_3651 : _GEN_280; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_282 = 8'h18 == auto_in_a_bits_source ? _T_3682 : _GEN_281; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_283 = 8'h19 == auto_in_a_bits_source ? _T_3713 : _GEN_282; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_284 = 8'h1a == auto_in_a_bits_source ? _T_3744 : _GEN_283; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_285 = 8'h1b == auto_in_a_bits_source ? _T_3775 : _GEN_284; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_286 = 8'h1c == auto_in_a_bits_source ? _T_3806 : _GEN_285; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_287 = 8'h1d == auto_in_a_bits_source ? _T_3837 : _GEN_286; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_288 = 8'h1e == auto_in_a_bits_source ? _T_3868 : _GEN_287; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_289 = 8'h1f == auto_in_a_bits_source ? _T_3899 : _GEN_288; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_290 = 8'h20 == auto_in_a_bits_source ? _T_3930 : _GEN_289; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_291 = 8'h21 == auto_in_a_bits_source ? _T_3961 : _GEN_290; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_292 = 8'h22 == auto_in_a_bits_source ? _T_3992 : _GEN_291; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_293 = 8'h23 == auto_in_a_bits_source ? _T_4023 : _GEN_292; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_294 = 8'h24 == auto_in_a_bits_source ? _T_4054 : _GEN_293; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_295 = 8'h25 == auto_in_a_bits_source ? _T_4085 : _GEN_294; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_296 = 8'h26 == auto_in_a_bits_source ? _T_4116 : _GEN_295; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_297 = 8'h27 == auto_in_a_bits_source ? _T_4147 : _GEN_296; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_298 = 8'h28 == auto_in_a_bits_source ? _T_4178 : _GEN_297; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_299 = 8'h29 == auto_in_a_bits_source ? _T_4209 : _GEN_298; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_300 = 8'h2a == auto_in_a_bits_source ? _T_4240 : _GEN_299; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_301 = 8'h2b == auto_in_a_bits_source ? _T_4271 : _GEN_300; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_302 = 8'h2c == auto_in_a_bits_source ? _T_4302 : _GEN_301; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_303 = 8'h2d == auto_in_a_bits_source ? _T_4333 : _GEN_302; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_304 = 8'h2e == auto_in_a_bits_source ? _T_4364 : _GEN_303; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_305 = 8'h2f == auto_in_a_bits_source ? _T_4395 : _GEN_304; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_306 = 8'h30 == auto_in_a_bits_source ? _T_4426 : _GEN_305; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_307 = 8'h31 == auto_in_a_bits_source ? _T_4457 : _GEN_306; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_308 = 8'h32 == auto_in_a_bits_source ? _T_4488 : _GEN_307; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_309 = 8'h33 == auto_in_a_bits_source ? _T_4519 : _GEN_308; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_310 = 8'h34 == auto_in_a_bits_source ? _T_4550 : _GEN_309; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_311 = 8'h35 == auto_in_a_bits_source ? _T_4581 : _GEN_310; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_312 = 8'h36 == auto_in_a_bits_source ? _T_4612 : _GEN_311; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_313 = 8'h37 == auto_in_a_bits_source ? _T_4643 : _GEN_312; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_314 = 8'h38 == auto_in_a_bits_source ? _T_4674 : _GEN_313; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_315 = 8'h39 == auto_in_a_bits_source ? _T_4705 : _GEN_314; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_316 = 8'h3a == auto_in_a_bits_source ? _T_4736 : _GEN_315; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_317 = 8'h3b == auto_in_a_bits_source ? _T_4767 : _GEN_316; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_318 = 8'h3c == auto_in_a_bits_source ? _T_4798 : _GEN_317; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_319 = 8'h3d == auto_in_a_bits_source ? _T_4829 : _GEN_318; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_320 = 8'h3e == auto_in_a_bits_source ? _T_4860 : _GEN_319; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_321 = 8'h3f == auto_in_a_bits_source ? _T_4891 : _GEN_320; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_322 = 8'h40 == auto_in_a_bits_source ? _T_4922 : _GEN_321; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_323 = 8'h41 == auto_in_a_bits_source ? _T_4953 : _GEN_322; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_324 = 8'h42 == auto_in_a_bits_source ? _T_4984 : _GEN_323; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_325 = 8'h43 == auto_in_a_bits_source ? _T_5015 : _GEN_324; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_326 = 8'h44 == auto_in_a_bits_source ? _T_5046 : _GEN_325; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_327 = 8'h45 == auto_in_a_bits_source ? _T_5077 : _GEN_326; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_328 = 8'h46 == auto_in_a_bits_source ? _T_5108 : _GEN_327; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_329 = 8'h47 == auto_in_a_bits_source ? _T_5139 : _GEN_328; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_330 = 8'h48 == auto_in_a_bits_source ? _T_5170 : _GEN_329; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_331 = 8'h49 == auto_in_a_bits_source ? _T_5201 : _GEN_330; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_332 = 8'h4a == auto_in_a_bits_source ? _T_5232 : _GEN_331; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_333 = 8'h4b == auto_in_a_bits_source ? _T_5263 : _GEN_332; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_334 = 8'h4c == auto_in_a_bits_source ? _T_5294 : _GEN_333; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_335 = 8'h4d == auto_in_a_bits_source ? _T_5325 : _GEN_334; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_336 = 8'h4e == auto_in_a_bits_source ? _T_5356 : _GEN_335; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_337 = 8'h4f == auto_in_a_bits_source ? _T_5387 : _GEN_336; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_338 = 8'h50 == auto_in_a_bits_source ? _T_5418 : _GEN_337; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_339 = 8'h51 == auto_in_a_bits_source ? _T_5449 : _GEN_338; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_340 = 8'h52 == auto_in_a_bits_source ? _T_5480 : _GEN_339; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_341 = 8'h53 == auto_in_a_bits_source ? _T_5511 : _GEN_340; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_342 = 8'h54 == auto_in_a_bits_source ? _T_5542 : _GEN_341; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_343 = 8'h55 == auto_in_a_bits_source ? _T_5573 : _GEN_342; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_344 = 8'h56 == auto_in_a_bits_source ? _T_5604 : _GEN_343; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_345 = 8'h57 == auto_in_a_bits_source ? _T_5635 : _GEN_344; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_346 = 8'h58 == auto_in_a_bits_source ? _T_5666 : _GEN_345; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_347 = 8'h59 == auto_in_a_bits_source ? _T_5697 : _GEN_346; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_348 = 8'h5a == auto_in_a_bits_source ? _T_5728 : _GEN_347; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_349 = 8'h5b == auto_in_a_bits_source ? _T_5759 : _GEN_348; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_350 = 8'h5c == auto_in_a_bits_source ? _T_5790 : _GEN_349; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_351 = 8'h5d == auto_in_a_bits_source ? _T_5821 : _GEN_350; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_352 = 8'h5e == auto_in_a_bits_source ? _T_5852 : _GEN_351; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_353 = 8'h5f == auto_in_a_bits_source ? _T_5883 : _GEN_352; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_354 = 8'h60 == auto_in_a_bits_source ? _T_5914 : _GEN_353; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_355 = 8'h61 == auto_in_a_bits_source ? _T_5945 : _GEN_354; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_356 = 8'h62 == auto_in_a_bits_source ? _T_5976 : _GEN_355; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_357 = 8'h63 == auto_in_a_bits_source ? _T_6007 : _GEN_356; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_358 = 8'h64 == auto_in_a_bits_source ? _T_6038 : _GEN_357; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_359 = 8'h65 == auto_in_a_bits_source ? _T_6069 : _GEN_358; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_360 = 8'h66 == auto_in_a_bits_source ? _T_6100 : _GEN_359; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_361 = 8'h67 == auto_in_a_bits_source ? _T_6131 : _GEN_360; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_362 = 8'h68 == auto_in_a_bits_source ? _T_6162 : _GEN_361; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_363 = 8'h69 == auto_in_a_bits_source ? _T_6193 : _GEN_362; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_364 = 8'h6a == auto_in_a_bits_source ? _T_6224 : _GEN_363; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_365 = 8'h6b == auto_in_a_bits_source ? _T_6255 : _GEN_364; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_366 = 8'h6c == auto_in_a_bits_source ? _T_6286 : _GEN_365; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_367 = 8'h6d == auto_in_a_bits_source ? _T_6317 : _GEN_366; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_368 = 8'h6e == auto_in_a_bits_source ? _T_6348 : _GEN_367; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_369 = 8'h6f == auto_in_a_bits_source ? _T_6379 : _GEN_368; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_370 = 8'h70 == auto_in_a_bits_source ? _T_6410 : _GEN_369; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_371 = 8'h71 == auto_in_a_bits_source ? _T_6441 : _GEN_370; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_372 = 8'h72 == auto_in_a_bits_source ? _T_6472 : _GEN_371; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_373 = 8'h73 == auto_in_a_bits_source ? _T_6503 : _GEN_372; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_374 = 8'h74 == auto_in_a_bits_source ? _T_6534 : _GEN_373; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_375 = 8'h75 == auto_in_a_bits_source ? _T_6565 : _GEN_374; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_376 = 8'h76 == auto_in_a_bits_source ? _T_6596 : _GEN_375; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_377 = 8'h77 == auto_in_a_bits_source ? _T_6627 : _GEN_376; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_378 = 8'h78 == auto_in_a_bits_source ? _T_6658 : _GEN_377; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_379 = 8'h79 == auto_in_a_bits_source ? _T_6689 : _GEN_378; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_380 = 8'h7a == auto_in_a_bits_source ? _T_6720 : _GEN_379; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_381 = 8'h7b == auto_in_a_bits_source ? _T_6751 : _GEN_380; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_382 = 8'h7c == auto_in_a_bits_source ? _T_6782 : _GEN_381; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_383 = 8'h7d == auto_in_a_bits_source ? _T_6813 : _GEN_382; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_384 = 8'h7e == auto_in_a_bits_source ? _T_6844 : _GEN_383; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_385 = 8'h7f == auto_in_a_bits_source ? _T_6875 : _GEN_384; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_386 = 8'h80 == auto_in_a_bits_source ? _T_6906 : _GEN_385; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_387 = 8'h81 == auto_in_a_bits_source ? _T_6937 : _GEN_386; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_388 = 8'h82 == auto_in_a_bits_source ? _T_6968 : _GEN_387; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_389 = 8'h83 == auto_in_a_bits_source ? _T_6999 : _GEN_388; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_390 = 8'h84 == auto_in_a_bits_source ? _T_7030 : _GEN_389; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_391 = 8'h85 == auto_in_a_bits_source ? _T_7061 : _GEN_390; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_392 = 8'h86 == auto_in_a_bits_source ? _T_7092 : _GEN_391; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_393 = 8'h87 == auto_in_a_bits_source ? _T_7123 : _GEN_392; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_394 = 8'h88 == auto_in_a_bits_source ? _T_7154 : _GEN_393; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_395 = 8'h89 == auto_in_a_bits_source ? _T_7185 : _GEN_394; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_396 = 8'h8a == auto_in_a_bits_source ? _T_7216 : _GEN_395; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_397 = 8'h8b == auto_in_a_bits_source ? _T_7247 : _GEN_396; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_398 = 8'h8c == auto_in_a_bits_source ? _T_7278 : _GEN_397; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_399 = 8'h8d == auto_in_a_bits_source ? _T_7309 : _GEN_398; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_400 = 8'h8e == auto_in_a_bits_source ? _T_7340 : _GEN_399; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_401 = 8'h8f == auto_in_a_bits_source ? _T_7371 : _GEN_400; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_402 = 8'h90 == auto_in_a_bits_source ? _T_7402 : _GEN_401; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_403 = 8'h91 == auto_in_a_bits_source ? _T_7433 : _GEN_402; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_404 = 8'h92 == auto_in_a_bits_source ? _T_7464 : _GEN_403; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_405 = 8'h93 == auto_in_a_bits_source ? _T_7495 : _GEN_404; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_406 = 8'h94 == auto_in_a_bits_source ? _T_7526 : _GEN_405; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_407 = 8'h95 == auto_in_a_bits_source ? _T_7557 : _GEN_406; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_408 = 8'h96 == auto_in_a_bits_source ? _T_7588 : _GEN_407; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_409 = 8'h97 == auto_in_a_bits_source ? _T_7619 : _GEN_408; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_410 = 8'h98 == auto_in_a_bits_source ? _T_7650 : _GEN_409; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_411 = 8'h99 == auto_in_a_bits_source ? _T_7681 : _GEN_410; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_412 = 8'h9a == auto_in_a_bits_source ? _T_7712 : _GEN_411; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_413 = 8'h9b == auto_in_a_bits_source ? _T_7743 : _GEN_412; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_414 = 8'h9c == auto_in_a_bits_source ? _T_7774 : _GEN_413; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_415 = 8'h9d == auto_in_a_bits_source ? _T_7805 : _GEN_414; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_416 = 8'h9e == auto_in_a_bits_source ? _T_7836 : _GEN_415; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_417 = 8'h9f == auto_in_a_bits_source ? _T_7867 : _GEN_416; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_418 = 8'ha0 == auto_in_a_bits_source ? _T_7898 : _GEN_417; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_419 = 8'ha1 == auto_in_a_bits_source ? _T_7929 : _GEN_418; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_420 = 8'ha2 == auto_in_a_bits_source ? _T_7960 : _GEN_419; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_421 = 8'ha3 == auto_in_a_bits_source ? _T_7991 : _GEN_420; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_422 = 8'ha4 == auto_in_a_bits_source ? _T_8022 : _GEN_421; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_423 = 8'ha5 == auto_in_a_bits_source ? _T_8053 : _GEN_422; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_424 = 8'ha6 == auto_in_a_bits_source ? _T_8084 : _GEN_423; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_425 = 8'ha7 == auto_in_a_bits_source ? _T_8115 : _GEN_424; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_426 = 8'ha8 == auto_in_a_bits_source ? _T_8146 : _GEN_425; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_427 = 8'ha9 == auto_in_a_bits_source ? _T_8177 : _GEN_426; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_428 = 8'haa == auto_in_a_bits_source ? _T_8208 : _GEN_427; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_429 = 8'hab == auto_in_a_bits_source ? _T_8239 : _GEN_428; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_430 = 8'hac == auto_in_a_bits_source ? _T_8270 : _GEN_429; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_431 = 8'had == auto_in_a_bits_source ? _T_8301 : _GEN_430; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_432 = 8'hae == auto_in_a_bits_source ? _T_8332 : _GEN_431; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_433 = 8'haf == auto_in_a_bits_source ? _T_8363 : _GEN_432; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_434 = 8'hb0 == auto_in_a_bits_source ? _T_8394 : _GEN_433; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_435 = 8'hb1 == auto_in_a_bits_source ? _T_8425 : _GEN_434; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_436 = 8'hb2 == auto_in_a_bits_source ? _T_8456 : _GEN_435; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_437 = 8'hb3 == auto_in_a_bits_source ? _T_8487 : _GEN_436; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_438 = 8'hb4 == auto_in_a_bits_source ? _T_8518 : _GEN_437; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_439 = 8'hb5 == auto_in_a_bits_source ? _T_8549 : _GEN_438; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_440 = 8'hb6 == auto_in_a_bits_source ? _T_8580 : _GEN_439; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_441 = 8'hb7 == auto_in_a_bits_source ? _T_8611 : _GEN_440; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_442 = 8'hb8 == auto_in_a_bits_source ? _T_8642 : _GEN_441; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_443 = 8'hb9 == auto_in_a_bits_source ? _T_8673 : _GEN_442; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_444 = 8'hba == auto_in_a_bits_source ? _T_8704 : _GEN_443; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_445 = 8'hbb == auto_in_a_bits_source ? _T_8735 : _GEN_444; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_446 = 8'hbc == auto_in_a_bits_source ? _T_8766 : _GEN_445; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_447 = 8'hbd == auto_in_a_bits_source ? _T_8797 : _GEN_446; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_448 = 8'hbe == auto_in_a_bits_source ? _T_8828 : _GEN_447; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_449 = 8'hbf == auto_in_a_bits_source ? _T_8859 : _GEN_448; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_450 = 8'hc0 == auto_in_a_bits_source ? _T_8890 : _GEN_449; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_451 = 8'hc1 == auto_in_a_bits_source ? _T_8921 : _GEN_450; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_452 = 8'hc2 == auto_in_a_bits_source ? _T_8952 : _GEN_451; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_453 = 8'hc3 == auto_in_a_bits_source ? _T_8983 : _GEN_452; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_454 = 8'hc4 == auto_in_a_bits_source ? _T_9014 : _GEN_453; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_455 = 8'hc5 == auto_in_a_bits_source ? _T_9045 : _GEN_454; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_456 = 8'hc6 == auto_in_a_bits_source ? _T_9076 : _GEN_455; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_457 = 8'hc7 == auto_in_a_bits_source ? _T_9107 : _GEN_456; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_458 = 8'hc8 == auto_in_a_bits_source ? _T_9138 : _GEN_457; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_459 = 8'hc9 == auto_in_a_bits_source ? _T_9169 : _GEN_458; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_460 = 8'hca == auto_in_a_bits_source ? _T_9200 : _GEN_459; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_461 = 8'hcb == auto_in_a_bits_source ? _T_9231 : _GEN_460; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_462 = 8'hcc == auto_in_a_bits_source ? _T_9262 : _GEN_461; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_463 = 8'hcd == auto_in_a_bits_source ? _T_9293 : _GEN_462; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_464 = 8'hce == auto_in_a_bits_source ? _T_9324 : _GEN_463; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_465 = 8'hcf == auto_in_a_bits_source ? _T_9355 : _GEN_464; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_466 = 8'hd0 == auto_in_a_bits_source ? _T_9386 : _GEN_465; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_467 = 8'hd1 == auto_in_a_bits_source ? _T_9417 : _GEN_466; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_468 = 8'hd2 == auto_in_a_bits_source ? _T_9448 : _GEN_467; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_469 = 8'hd3 == auto_in_a_bits_source ? _T_9479 : _GEN_468; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_470 = 8'hd4 == auto_in_a_bits_source ? _T_9510 : _GEN_469; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_471 = 8'hd5 == auto_in_a_bits_source ? _T_9541 : _GEN_470; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_472 = 8'hd6 == auto_in_a_bits_source ? _T_9572 : _GEN_471; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_473 = 8'hd7 == auto_in_a_bits_source ? _T_9603 : _GEN_472; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_474 = 8'hd8 == auto_in_a_bits_source ? _T_9634 : _GEN_473; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_475 = 8'hd9 == auto_in_a_bits_source ? _T_9665 : _GEN_474; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_476 = 8'hda == auto_in_a_bits_source ? _T_9696 : _GEN_475; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_477 = 8'hdb == auto_in_a_bits_source ? _T_9727 : _GEN_476; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_478 = 8'hdc == auto_in_a_bits_source ? _T_9758 : _GEN_477; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_479 = 8'hdd == auto_in_a_bits_source ? _T_9789 : _GEN_478; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_480 = 8'hde == auto_in_a_bits_source ? _T_9820 : _GEN_479; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_481 = 8'hdf == auto_in_a_bits_source ? _T_9851 : _GEN_480; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_482 = 8'he0 == auto_in_a_bits_source ? _T_9882 : _GEN_481; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_483 = 8'he1 == auto_in_a_bits_source ? _T_9913 : _GEN_482; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_484 = 8'he2 == auto_in_a_bits_source ? _T_9944 : _GEN_483; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_485 = 8'he3 == auto_in_a_bits_source ? _T_9975 : _GEN_484; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_486 = 8'he4 == auto_in_a_bits_source ? _T_10006 : _GEN_485; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_487 = 8'he5 == auto_in_a_bits_source ? _T_10037 : _GEN_486; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_488 = 8'he6 == auto_in_a_bits_source ? _T_10068 : _GEN_487; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_489 = 8'he7 == auto_in_a_bits_source ? _T_10099 : _GEN_488; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_490 = 8'he8 == auto_in_a_bits_source ? _T_10130 : _GEN_489; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_491 = 8'he9 == auto_in_a_bits_source ? _T_10161 : _GEN_490; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_492 = 8'hea == auto_in_a_bits_source ? _T_10192 : _GEN_491; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_493 = 8'heb == auto_in_a_bits_source ? _T_10223 : _GEN_492; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_494 = 8'hec == auto_in_a_bits_source ? _T_10254 : _GEN_493; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_495 = 8'hed == auto_in_a_bits_source ? _T_10285 : _GEN_494; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_496 = 8'hee == auto_in_a_bits_source ? _T_10316 : _GEN_495; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_497 = 8'hef == auto_in_a_bits_source ? _T_10347 : _GEN_496; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_498 = 8'hf0 == auto_in_a_bits_source ? _T_10378 : _GEN_497; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_499 = 8'hf1 == auto_in_a_bits_source ? _T_10409 : _GEN_498; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_500 = 8'hf2 == auto_in_a_bits_source ? _T_10440 : _GEN_499; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_501 = 8'hf3 == auto_in_a_bits_source ? _T_10471 : _GEN_500; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_502 = 8'hf4 == auto_in_a_bits_source ? _T_10502 : _GEN_501; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_503 = 8'hf5 == auto_in_a_bits_source ? _T_10533 : _GEN_502; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_504 = 8'hf6 == auto_in_a_bits_source ? _T_10564 : _GEN_503; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_505 = 8'hf7 == auto_in_a_bits_source ? _T_10595 : _GEN_504; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_506 = 8'hf8 == auto_in_a_bits_source ? _T_10626 : _GEN_505; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_507 = 8'hf9 == auto_in_a_bits_source ? _T_10657 : _GEN_506; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_508 = 8'hfa == auto_in_a_bits_source ? _T_10688 : _GEN_507; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_509 = 8'hfb == auto_in_a_bits_source ? _T_10719 : _GEN_508; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_510 = 8'hfc == auto_in_a_bits_source ? _T_10750 : _GEN_509; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_511 = 8'hfd == auto_in_a_bits_source ? _T_10781 : _GEN_510; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_512 = 8'hfe == auto_in_a_bits_source ? _T_10812 : _GEN_511; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _GEN_513 = 8'hff == auto_in_a_bits_source ? _T_10843 : _GEN_512; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _T_2311 = _T_2307 == 3'h0; // @[Edges.scala 231:25:boom.system.TestHarness.MegaBoomConfig.fir@20247.4]
  assign _T_2377 = _GEN_513 & _T_2311; // @[ToAXI4.scala 176:49:boom.system.TestHarness.MegaBoomConfig.fir@20363.4]
  assign _T_2378 = _T_2377 == 1'h0; // @[ToAXI4.scala 177:21:boom.system.TestHarness.MegaBoomConfig.fir@20364.4]
  assign _T_2338_ready = Queue_1_io_enq_ready; // @[ToAXI4.scala 146:25:boom.system.TestHarness.MegaBoomConfig.fir@20281.4 Decoupled.scala 296:17:boom.system.TestHarness.MegaBoomConfig.fir@20315.4]
  assign _T_2379 = _T_2365 | _T_2338_ready; // @[ToAXI4.scala 177:52:boom.system.TestHarness.MegaBoomConfig.fir@20365.4]
  assign _T_2341_ready = Queue_io_enq_ready; // @[ToAXI4.scala 147:23:boom.system.TestHarness.MegaBoomConfig.fir@20283.4 Decoupled.scala 296:17:boom.system.TestHarness.MegaBoomConfig.fir@20292.4]
  assign _T_2380 = _T_2379 & _T_2341_ready; // @[ToAXI4.scala 177:70:boom.system.TestHarness.MegaBoomConfig.fir@20366.4]
  assign _T_2381 = _T_2296 ? _T_2380 : _T_2338_ready; // @[ToAXI4.scala 177:34:boom.system.TestHarness.MegaBoomConfig.fir@20367.4]
  assign _T_2382 = _T_2378 & _T_2381; // @[ToAXI4.scala 177:28:boom.system.TestHarness.MegaBoomConfig.fir@20368.4]
  assign _T_2297 = _T_2382 & auto_in_a_valid; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@20234.4]
  assign _T_2299 = 13'h3f << auto_in_a_bits_size; // @[package.scala 185:77:boom.system.TestHarness.MegaBoomConfig.fir@20236.4]
  assign _T_2300 = _T_2299[5:0]; // @[package.scala 185:82:boom.system.TestHarness.MegaBoomConfig.fir@20237.4]
  assign _T_2301 = ~ _T_2300; // @[package.scala 185:46:boom.system.TestHarness.MegaBoomConfig.fir@20238.4]
  assign _T_2302 = _T_2301[5:3]; // @[Edges.scala 220:59:boom.system.TestHarness.MegaBoomConfig.fir@20239.4]
  assign _T_2305 = _T_2296 ? _T_2302 : 3'h0; // @[Edges.scala 221:14:boom.system.TestHarness.MegaBoomConfig.fir@20242.4]
  assign _T_2308 = _T_2307 - 3'h1; // @[Edges.scala 230:28:boom.system.TestHarness.MegaBoomConfig.fir@20244.4]
  assign _T_2309 = $unsigned(_T_2308); // @[Edges.scala 230:28:boom.system.TestHarness.MegaBoomConfig.fir@20245.4]
  assign _T_2310 = _T_2309[2:0]; // @[Edges.scala 230:28:boom.system.TestHarness.MegaBoomConfig.fir@20246.4]
  assign _T_2312 = _T_2307 == 3'h1; // @[Edges.scala 232:25:boom.system.TestHarness.MegaBoomConfig.fir@20248.4]
  assign _T_2313 = _T_2305 == 3'h0; // @[Edges.scala 232:47:boom.system.TestHarness.MegaBoomConfig.fir@20249.4]
  assign _T_2314 = _T_2312 | _T_2313; // @[Edges.scala 232:37:boom.system.TestHarness.MegaBoomConfig.fir@20250.4]
  assign _GEN_773 = {{8'd0}, auto_in_a_bits_size}; // @[ToAXI4.scala 134:55:boom.system.TestHarness.MegaBoomConfig.fir@20275.4]
  assign _T_2328 = _GEN_773 << 8; // @[ToAXI4.scala 134:55:boom.system.TestHarness.MegaBoomConfig.fir@20275.4]
  assign _GEN_774 = {{3'd0}, auto_in_a_bits_source}; // @[ToAXI4.scala 134:45:boom.system.TestHarness.MegaBoomConfig.fir@20276.4]
  assign _T_2329 = _GEN_774 | _T_2328; // @[ToAXI4.scala 134:45:boom.system.TestHarness.MegaBoomConfig.fir@20276.4]
  assign _T_2330 = auto_out_r_bits_user[7:0]; // @[ToAXI4.scala 137:50:boom.system.TestHarness.MegaBoomConfig.fir@20277.4]
  assign _T_2331 = auto_out_r_bits_user[10:8]; // @[ToAXI4.scala 138:50:boom.system.TestHarness.MegaBoomConfig.fir@20278.4]
  assign _T_2332 = auto_out_b_bits_user[7:0]; // @[ToAXI4.scala 141:50:boom.system.TestHarness.MegaBoomConfig.fir@20279.4]
  assign _T_2333 = auto_out_b_bits_user[10:8]; // @[ToAXI4.scala 142:50:boom.system.TestHarness.MegaBoomConfig.fir@20280.4]
  assign _T_2356_bits_wen = Queue_1_io_deq_bits_wen; // @[Decoupled.scala 314:19:boom.system.TestHarness.MegaBoomConfig.fir@20316.4 Decoupled.scala 315:14:boom.system.TestHarness.MegaBoomConfig.fir@20317.4]
  assign _T_2360 = _T_2356_bits_wen == 1'h0; // @[ToAXI4.scala 154:42:boom.system.TestHarness.MegaBoomConfig.fir@20332.4]
  assign _T_2356_valid = Queue_1_io_deq_valid; // @[Decoupled.scala 314:19:boom.system.TestHarness.MegaBoomConfig.fir@20316.4 Decoupled.scala 316:15:boom.system.TestHarness.MegaBoomConfig.fir@20328.4]
  assign _T_2367 = _T_2314 == 1'h0; // @[ToAXI4.scala 161:38:boom.system.TestHarness.MegaBoomConfig.fir@20342.6]
  assign _GEN_3 = 8'h1 == auto_in_a_bits_source ? 8'h1 : 8'h0; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_4 = 8'h2 == auto_in_a_bits_source ? 8'h2 : _GEN_3; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_5 = 8'h3 == auto_in_a_bits_source ? 8'h3 : _GEN_4; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_6 = 8'h4 == auto_in_a_bits_source ? 8'h4 : _GEN_5; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_7 = 8'h5 == auto_in_a_bits_source ? 8'h5 : _GEN_6; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_8 = 8'h6 == auto_in_a_bits_source ? 8'h6 : _GEN_7; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_9 = 8'h7 == auto_in_a_bits_source ? 8'h7 : _GEN_8; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_10 = 8'h8 == auto_in_a_bits_source ? 8'h8 : _GEN_9; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_11 = 8'h9 == auto_in_a_bits_source ? 8'h9 : _GEN_10; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_12 = 8'ha == auto_in_a_bits_source ? 8'ha : _GEN_11; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_13 = 8'hb == auto_in_a_bits_source ? 8'hb : _GEN_12; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_14 = 8'hc == auto_in_a_bits_source ? 8'hc : _GEN_13; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_15 = 8'hd == auto_in_a_bits_source ? 8'hd : _GEN_14; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_16 = 8'he == auto_in_a_bits_source ? 8'he : _GEN_15; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_17 = 8'hf == auto_in_a_bits_source ? 8'hf : _GEN_16; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_18 = 8'h10 == auto_in_a_bits_source ? 8'h10 : _GEN_17; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_19 = 8'h11 == auto_in_a_bits_source ? 8'h11 : _GEN_18; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_20 = 8'h12 == auto_in_a_bits_source ? 8'h12 : _GEN_19; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_21 = 8'h13 == auto_in_a_bits_source ? 8'h13 : _GEN_20; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_22 = 8'h14 == auto_in_a_bits_source ? 8'h14 : _GEN_21; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_23 = 8'h15 == auto_in_a_bits_source ? 8'h15 : _GEN_22; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_24 = 8'h16 == auto_in_a_bits_source ? 8'h16 : _GEN_23; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_25 = 8'h17 == auto_in_a_bits_source ? 8'h17 : _GEN_24; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_26 = 8'h18 == auto_in_a_bits_source ? 8'h18 : _GEN_25; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_27 = 8'h19 == auto_in_a_bits_source ? 8'h19 : _GEN_26; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_28 = 8'h1a == auto_in_a_bits_source ? 8'h1a : _GEN_27; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_29 = 8'h1b == auto_in_a_bits_source ? 8'h1b : _GEN_28; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_30 = 8'h1c == auto_in_a_bits_source ? 8'h1c : _GEN_29; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_31 = 8'h1d == auto_in_a_bits_source ? 8'h1d : _GEN_30; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_32 = 8'h1e == auto_in_a_bits_source ? 8'h1e : _GEN_31; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_33 = 8'h1f == auto_in_a_bits_source ? 8'h1f : _GEN_32; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_34 = 8'h20 == auto_in_a_bits_source ? 8'h20 : _GEN_33; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_35 = 8'h21 == auto_in_a_bits_source ? 8'h21 : _GEN_34; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_36 = 8'h22 == auto_in_a_bits_source ? 8'h22 : _GEN_35; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_37 = 8'h23 == auto_in_a_bits_source ? 8'h23 : _GEN_36; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_38 = 8'h24 == auto_in_a_bits_source ? 8'h24 : _GEN_37; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_39 = 8'h25 == auto_in_a_bits_source ? 8'h25 : _GEN_38; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_40 = 8'h26 == auto_in_a_bits_source ? 8'h26 : _GEN_39; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_41 = 8'h27 == auto_in_a_bits_source ? 8'h27 : _GEN_40; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_42 = 8'h28 == auto_in_a_bits_source ? 8'h28 : _GEN_41; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_43 = 8'h29 == auto_in_a_bits_source ? 8'h29 : _GEN_42; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_44 = 8'h2a == auto_in_a_bits_source ? 8'h2a : _GEN_43; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_45 = 8'h2b == auto_in_a_bits_source ? 8'h2b : _GEN_44; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_46 = 8'h2c == auto_in_a_bits_source ? 8'h2c : _GEN_45; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_47 = 8'h2d == auto_in_a_bits_source ? 8'h2d : _GEN_46; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_48 = 8'h2e == auto_in_a_bits_source ? 8'h2e : _GEN_47; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_49 = 8'h2f == auto_in_a_bits_source ? 8'h2f : _GEN_48; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_50 = 8'h30 == auto_in_a_bits_source ? 8'h30 : _GEN_49; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_51 = 8'h31 == auto_in_a_bits_source ? 8'h31 : _GEN_50; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_52 = 8'h32 == auto_in_a_bits_source ? 8'h32 : _GEN_51; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_53 = 8'h33 == auto_in_a_bits_source ? 8'h33 : _GEN_52; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_54 = 8'h34 == auto_in_a_bits_source ? 8'h34 : _GEN_53; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_55 = 8'h35 == auto_in_a_bits_source ? 8'h35 : _GEN_54; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_56 = 8'h36 == auto_in_a_bits_source ? 8'h36 : _GEN_55; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_57 = 8'h37 == auto_in_a_bits_source ? 8'h37 : _GEN_56; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_58 = 8'h38 == auto_in_a_bits_source ? 8'h38 : _GEN_57; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_59 = 8'h39 == auto_in_a_bits_source ? 8'h39 : _GEN_58; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_60 = 8'h3a == auto_in_a_bits_source ? 8'h3a : _GEN_59; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_61 = 8'h3b == auto_in_a_bits_source ? 8'h3b : _GEN_60; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_62 = 8'h3c == auto_in_a_bits_source ? 8'h3c : _GEN_61; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_63 = 8'h3d == auto_in_a_bits_source ? 8'h3d : _GEN_62; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_64 = 8'h3e == auto_in_a_bits_source ? 8'h3e : _GEN_63; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_65 = 8'h3f == auto_in_a_bits_source ? 8'h3f : _GEN_64; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_66 = 8'h40 == auto_in_a_bits_source ? 8'h40 : _GEN_65; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_67 = 8'h41 == auto_in_a_bits_source ? 8'h41 : _GEN_66; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_68 = 8'h42 == auto_in_a_bits_source ? 8'h42 : _GEN_67; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_69 = 8'h43 == auto_in_a_bits_source ? 8'h43 : _GEN_68; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_70 = 8'h44 == auto_in_a_bits_source ? 8'h44 : _GEN_69; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_71 = 8'h45 == auto_in_a_bits_source ? 8'h45 : _GEN_70; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_72 = 8'h46 == auto_in_a_bits_source ? 8'h46 : _GEN_71; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_73 = 8'h47 == auto_in_a_bits_source ? 8'h47 : _GEN_72; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_74 = 8'h48 == auto_in_a_bits_source ? 8'h48 : _GEN_73; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_75 = 8'h49 == auto_in_a_bits_source ? 8'h49 : _GEN_74; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_76 = 8'h4a == auto_in_a_bits_source ? 8'h4a : _GEN_75; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_77 = 8'h4b == auto_in_a_bits_source ? 8'h4b : _GEN_76; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_78 = 8'h4c == auto_in_a_bits_source ? 8'h4c : _GEN_77; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_79 = 8'h4d == auto_in_a_bits_source ? 8'h4d : _GEN_78; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_80 = 8'h4e == auto_in_a_bits_source ? 8'h4e : _GEN_79; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_81 = 8'h4f == auto_in_a_bits_source ? 8'h4f : _GEN_80; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_82 = 8'h50 == auto_in_a_bits_source ? 8'h50 : _GEN_81; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_83 = 8'h51 == auto_in_a_bits_source ? 8'h51 : _GEN_82; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_84 = 8'h52 == auto_in_a_bits_source ? 8'h52 : _GEN_83; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_85 = 8'h53 == auto_in_a_bits_source ? 8'h53 : _GEN_84; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_86 = 8'h54 == auto_in_a_bits_source ? 8'h54 : _GEN_85; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_87 = 8'h55 == auto_in_a_bits_source ? 8'h55 : _GEN_86; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_88 = 8'h56 == auto_in_a_bits_source ? 8'h56 : _GEN_87; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_89 = 8'h57 == auto_in_a_bits_source ? 8'h57 : _GEN_88; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_90 = 8'h58 == auto_in_a_bits_source ? 8'h58 : _GEN_89; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_91 = 8'h59 == auto_in_a_bits_source ? 8'h59 : _GEN_90; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_92 = 8'h5a == auto_in_a_bits_source ? 8'h5a : _GEN_91; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_93 = 8'h5b == auto_in_a_bits_source ? 8'h5b : _GEN_92; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_94 = 8'h5c == auto_in_a_bits_source ? 8'h5c : _GEN_93; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_95 = 8'h5d == auto_in_a_bits_source ? 8'h5d : _GEN_94; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_96 = 8'h5e == auto_in_a_bits_source ? 8'h5e : _GEN_95; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_97 = 8'h5f == auto_in_a_bits_source ? 8'h5f : _GEN_96; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_98 = 8'h60 == auto_in_a_bits_source ? 8'h60 : _GEN_97; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_99 = 8'h61 == auto_in_a_bits_source ? 8'h61 : _GEN_98; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_100 = 8'h62 == auto_in_a_bits_source ? 8'h62 : _GEN_99; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_101 = 8'h63 == auto_in_a_bits_source ? 8'h63 : _GEN_100; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_102 = 8'h64 == auto_in_a_bits_source ? 8'h64 : _GEN_101; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_103 = 8'h65 == auto_in_a_bits_source ? 8'h65 : _GEN_102; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_104 = 8'h66 == auto_in_a_bits_source ? 8'h66 : _GEN_103; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_105 = 8'h67 == auto_in_a_bits_source ? 8'h67 : _GEN_104; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_106 = 8'h68 == auto_in_a_bits_source ? 8'h68 : _GEN_105; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_107 = 8'h69 == auto_in_a_bits_source ? 8'h69 : _GEN_106; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_108 = 8'h6a == auto_in_a_bits_source ? 8'h6a : _GEN_107; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_109 = 8'h6b == auto_in_a_bits_source ? 8'h6b : _GEN_108; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_110 = 8'h6c == auto_in_a_bits_source ? 8'h6c : _GEN_109; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_111 = 8'h6d == auto_in_a_bits_source ? 8'h6d : _GEN_110; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_112 = 8'h6e == auto_in_a_bits_source ? 8'h6e : _GEN_111; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_113 = 8'h6f == auto_in_a_bits_source ? 8'h6f : _GEN_112; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_114 = 8'h70 == auto_in_a_bits_source ? 8'h70 : _GEN_113; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_115 = 8'h71 == auto_in_a_bits_source ? 8'h71 : _GEN_114; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_116 = 8'h72 == auto_in_a_bits_source ? 8'h72 : _GEN_115; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_117 = 8'h73 == auto_in_a_bits_source ? 8'h73 : _GEN_116; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_118 = 8'h74 == auto_in_a_bits_source ? 8'h74 : _GEN_117; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_119 = 8'h75 == auto_in_a_bits_source ? 8'h75 : _GEN_118; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_120 = 8'h76 == auto_in_a_bits_source ? 8'h76 : _GEN_119; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_121 = 8'h77 == auto_in_a_bits_source ? 8'h77 : _GEN_120; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_122 = 8'h78 == auto_in_a_bits_source ? 8'h78 : _GEN_121; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_123 = 8'h79 == auto_in_a_bits_source ? 8'h79 : _GEN_122; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_124 = 8'h7a == auto_in_a_bits_source ? 8'h7a : _GEN_123; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_125 = 8'h7b == auto_in_a_bits_source ? 8'h7b : _GEN_124; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_126 = 8'h7c == auto_in_a_bits_source ? 8'h7c : _GEN_125; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_127 = 8'h7d == auto_in_a_bits_source ? 8'h7d : _GEN_126; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_128 = 8'h7e == auto_in_a_bits_source ? 8'h7e : _GEN_127; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_129 = 8'h7f == auto_in_a_bits_source ? 8'h7f : _GEN_128; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_130 = 8'h80 == auto_in_a_bits_source ? 8'h80 : _GEN_129; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_131 = 8'h81 == auto_in_a_bits_source ? 8'h81 : _GEN_130; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_132 = 8'h82 == auto_in_a_bits_source ? 8'h82 : _GEN_131; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_133 = 8'h83 == auto_in_a_bits_source ? 8'h83 : _GEN_132; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_134 = 8'h84 == auto_in_a_bits_source ? 8'h84 : _GEN_133; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_135 = 8'h85 == auto_in_a_bits_source ? 8'h85 : _GEN_134; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_136 = 8'h86 == auto_in_a_bits_source ? 8'h86 : _GEN_135; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_137 = 8'h87 == auto_in_a_bits_source ? 8'h87 : _GEN_136; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_138 = 8'h88 == auto_in_a_bits_source ? 8'h88 : _GEN_137; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_139 = 8'h89 == auto_in_a_bits_source ? 8'h89 : _GEN_138; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_140 = 8'h8a == auto_in_a_bits_source ? 8'h8a : _GEN_139; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_141 = 8'h8b == auto_in_a_bits_source ? 8'h8b : _GEN_140; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_142 = 8'h8c == auto_in_a_bits_source ? 8'h8c : _GEN_141; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_143 = 8'h8d == auto_in_a_bits_source ? 8'h8d : _GEN_142; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_144 = 8'h8e == auto_in_a_bits_source ? 8'h8e : _GEN_143; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_145 = 8'h8f == auto_in_a_bits_source ? 8'h8f : _GEN_144; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_146 = 8'h90 == auto_in_a_bits_source ? 8'h90 : _GEN_145; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_147 = 8'h91 == auto_in_a_bits_source ? 8'h91 : _GEN_146; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_148 = 8'h92 == auto_in_a_bits_source ? 8'h92 : _GEN_147; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_149 = 8'h93 == auto_in_a_bits_source ? 8'h93 : _GEN_148; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_150 = 8'h94 == auto_in_a_bits_source ? 8'h94 : _GEN_149; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_151 = 8'h95 == auto_in_a_bits_source ? 8'h95 : _GEN_150; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_152 = 8'h96 == auto_in_a_bits_source ? 8'h96 : _GEN_151; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_153 = 8'h97 == auto_in_a_bits_source ? 8'h97 : _GEN_152; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_154 = 8'h98 == auto_in_a_bits_source ? 8'h98 : _GEN_153; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_155 = 8'h99 == auto_in_a_bits_source ? 8'h99 : _GEN_154; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_156 = 8'h9a == auto_in_a_bits_source ? 8'h9a : _GEN_155; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_157 = 8'h9b == auto_in_a_bits_source ? 8'h9b : _GEN_156; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_158 = 8'h9c == auto_in_a_bits_source ? 8'h9c : _GEN_157; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_159 = 8'h9d == auto_in_a_bits_source ? 8'h9d : _GEN_158; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_160 = 8'h9e == auto_in_a_bits_source ? 8'h9e : _GEN_159; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_161 = 8'h9f == auto_in_a_bits_source ? 8'h9f : _GEN_160; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_162 = 8'ha0 == auto_in_a_bits_source ? 8'ha0 : _GEN_161; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_163 = 8'ha1 == auto_in_a_bits_source ? 8'ha1 : _GEN_162; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_164 = 8'ha2 == auto_in_a_bits_source ? 8'ha2 : _GEN_163; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_165 = 8'ha3 == auto_in_a_bits_source ? 8'ha3 : _GEN_164; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_166 = 8'ha4 == auto_in_a_bits_source ? 8'ha4 : _GEN_165; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_167 = 8'ha5 == auto_in_a_bits_source ? 8'ha5 : _GEN_166; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_168 = 8'ha6 == auto_in_a_bits_source ? 8'ha6 : _GEN_167; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_169 = 8'ha7 == auto_in_a_bits_source ? 8'ha7 : _GEN_168; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_170 = 8'ha8 == auto_in_a_bits_source ? 8'ha8 : _GEN_169; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_171 = 8'ha9 == auto_in_a_bits_source ? 8'ha9 : _GEN_170; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_172 = 8'haa == auto_in_a_bits_source ? 8'haa : _GEN_171; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_173 = 8'hab == auto_in_a_bits_source ? 8'hab : _GEN_172; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_174 = 8'hac == auto_in_a_bits_source ? 8'hac : _GEN_173; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_175 = 8'had == auto_in_a_bits_source ? 8'had : _GEN_174; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_176 = 8'hae == auto_in_a_bits_source ? 8'hae : _GEN_175; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_177 = 8'haf == auto_in_a_bits_source ? 8'haf : _GEN_176; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_178 = 8'hb0 == auto_in_a_bits_source ? 8'hb0 : _GEN_177; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_179 = 8'hb1 == auto_in_a_bits_source ? 8'hb1 : _GEN_178; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_180 = 8'hb2 == auto_in_a_bits_source ? 8'hb2 : _GEN_179; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_181 = 8'hb3 == auto_in_a_bits_source ? 8'hb3 : _GEN_180; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_182 = 8'hb4 == auto_in_a_bits_source ? 8'hb4 : _GEN_181; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_183 = 8'hb5 == auto_in_a_bits_source ? 8'hb5 : _GEN_182; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_184 = 8'hb6 == auto_in_a_bits_source ? 8'hb6 : _GEN_183; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_185 = 8'hb7 == auto_in_a_bits_source ? 8'hb7 : _GEN_184; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_186 = 8'hb8 == auto_in_a_bits_source ? 8'hb8 : _GEN_185; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_187 = 8'hb9 == auto_in_a_bits_source ? 8'hb9 : _GEN_186; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_188 = 8'hba == auto_in_a_bits_source ? 8'hba : _GEN_187; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_189 = 8'hbb == auto_in_a_bits_source ? 8'hbb : _GEN_188; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_190 = 8'hbc == auto_in_a_bits_source ? 8'hbc : _GEN_189; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_191 = 8'hbd == auto_in_a_bits_source ? 8'hbd : _GEN_190; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_192 = 8'hbe == auto_in_a_bits_source ? 8'hbe : _GEN_191; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_193 = 8'hbf == auto_in_a_bits_source ? 8'hbf : _GEN_192; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_194 = 8'hc0 == auto_in_a_bits_source ? 8'hc0 : _GEN_193; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_195 = 8'hc1 == auto_in_a_bits_source ? 8'hc1 : _GEN_194; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_196 = 8'hc2 == auto_in_a_bits_source ? 8'hc2 : _GEN_195; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_197 = 8'hc3 == auto_in_a_bits_source ? 8'hc3 : _GEN_196; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_198 = 8'hc4 == auto_in_a_bits_source ? 8'hc4 : _GEN_197; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_199 = 8'hc5 == auto_in_a_bits_source ? 8'hc5 : _GEN_198; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_200 = 8'hc6 == auto_in_a_bits_source ? 8'hc6 : _GEN_199; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_201 = 8'hc7 == auto_in_a_bits_source ? 8'hc7 : _GEN_200; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_202 = 8'hc8 == auto_in_a_bits_source ? 8'hc8 : _GEN_201; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_203 = 8'hc9 == auto_in_a_bits_source ? 8'hc9 : _GEN_202; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_204 = 8'hca == auto_in_a_bits_source ? 8'hca : _GEN_203; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_205 = 8'hcb == auto_in_a_bits_source ? 8'hcb : _GEN_204; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_206 = 8'hcc == auto_in_a_bits_source ? 8'hcc : _GEN_205; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_207 = 8'hcd == auto_in_a_bits_source ? 8'hcd : _GEN_206; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_208 = 8'hce == auto_in_a_bits_source ? 8'hce : _GEN_207; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_209 = 8'hcf == auto_in_a_bits_source ? 8'hcf : _GEN_208; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_210 = 8'hd0 == auto_in_a_bits_source ? 8'hd0 : _GEN_209; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_211 = 8'hd1 == auto_in_a_bits_source ? 8'hd1 : _GEN_210; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_212 = 8'hd2 == auto_in_a_bits_source ? 8'hd2 : _GEN_211; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_213 = 8'hd3 == auto_in_a_bits_source ? 8'hd3 : _GEN_212; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_214 = 8'hd4 == auto_in_a_bits_source ? 8'hd4 : _GEN_213; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_215 = 8'hd5 == auto_in_a_bits_source ? 8'hd5 : _GEN_214; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_216 = 8'hd6 == auto_in_a_bits_source ? 8'hd6 : _GEN_215; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_217 = 8'hd7 == auto_in_a_bits_source ? 8'hd7 : _GEN_216; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_218 = 8'hd8 == auto_in_a_bits_source ? 8'hd8 : _GEN_217; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_219 = 8'hd9 == auto_in_a_bits_source ? 8'hd9 : _GEN_218; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_220 = 8'hda == auto_in_a_bits_source ? 8'hda : _GEN_219; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_221 = 8'hdb == auto_in_a_bits_source ? 8'hdb : _GEN_220; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_222 = 8'hdc == auto_in_a_bits_source ? 8'hdc : _GEN_221; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_223 = 8'hdd == auto_in_a_bits_source ? 8'hdd : _GEN_222; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_224 = 8'hde == auto_in_a_bits_source ? 8'hde : _GEN_223; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_225 = 8'hdf == auto_in_a_bits_source ? 8'hdf : _GEN_224; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_226 = 8'he0 == auto_in_a_bits_source ? 8'he0 : _GEN_225; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_227 = 8'he1 == auto_in_a_bits_source ? 8'he1 : _GEN_226; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_228 = 8'he2 == auto_in_a_bits_source ? 8'he2 : _GEN_227; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_229 = 8'he3 == auto_in_a_bits_source ? 8'he3 : _GEN_228; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_230 = 8'he4 == auto_in_a_bits_source ? 8'he4 : _GEN_229; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_231 = 8'he5 == auto_in_a_bits_source ? 8'he5 : _GEN_230; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_232 = 8'he6 == auto_in_a_bits_source ? 8'he6 : _GEN_231; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_233 = 8'he7 == auto_in_a_bits_source ? 8'he7 : _GEN_232; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_234 = 8'he8 == auto_in_a_bits_source ? 8'he8 : _GEN_233; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_235 = 8'he9 == auto_in_a_bits_source ? 8'he9 : _GEN_234; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_236 = 8'hea == auto_in_a_bits_source ? 8'hea : _GEN_235; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_237 = 8'heb == auto_in_a_bits_source ? 8'heb : _GEN_236; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_238 = 8'hec == auto_in_a_bits_source ? 8'hec : _GEN_237; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_239 = 8'hed == auto_in_a_bits_source ? 8'hed : _GEN_238; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_240 = 8'hee == auto_in_a_bits_source ? 8'hee : _GEN_239; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_241 = 8'hef == auto_in_a_bits_source ? 8'hef : _GEN_240; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_242 = 8'hf0 == auto_in_a_bits_source ? 8'hf0 : _GEN_241; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_243 = 8'hf1 == auto_in_a_bits_source ? 8'hf1 : _GEN_242; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_244 = 8'hf2 == auto_in_a_bits_source ? 8'hf2 : _GEN_243; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_245 = 8'hf3 == auto_in_a_bits_source ? 8'hf3 : _GEN_244; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_246 = 8'hf4 == auto_in_a_bits_source ? 8'hf4 : _GEN_245; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_247 = 8'hf5 == auto_in_a_bits_source ? 8'hf5 : _GEN_246; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_248 = 8'hf6 == auto_in_a_bits_source ? 8'hf6 : _GEN_247; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_249 = 8'hf7 == auto_in_a_bits_source ? 8'hf7 : _GEN_248; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_250 = 8'hf8 == auto_in_a_bits_source ? 8'hf8 : _GEN_249; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_251 = 8'hf9 == auto_in_a_bits_source ? 8'hf9 : _GEN_250; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_252 = 8'hfa == auto_in_a_bits_source ? 8'hfa : _GEN_251; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_253 = 8'hfb == auto_in_a_bits_source ? 8'hfb : _GEN_252; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_254 = 8'hfc == auto_in_a_bits_source ? 8'hfc : _GEN_253; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_255 = 8'hfd == auto_in_a_bits_source ? 8'hfd : _GEN_254; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_256 = 8'hfe == auto_in_a_bits_source ? 8'hfe : _GEN_255; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _GEN_257 = 8'hff == auto_in_a_bits_source ? 8'hff : _GEN_256; // @[ToAXI4.scala 165:17:boom.system.TestHarness.MegaBoomConfig.fir@20346.4]
  assign _T_2370 = 18'h7ff << auto_in_a_bits_size; // @[package.scala 185:77:boom.system.TestHarness.MegaBoomConfig.fir@20349.4]
  assign _T_2371 = _T_2370[10:0]; // @[package.scala 185:82:boom.system.TestHarness.MegaBoomConfig.fir@20350.4]
  assign _T_2372 = ~ _T_2371; // @[package.scala 185:46:boom.system.TestHarness.MegaBoomConfig.fir@20351.4]
  assign _T_2374 = auto_in_a_bits_size >= 3'h3; // @[ToAXI4.scala 168:31:boom.system.TestHarness.MegaBoomConfig.fir@20354.4]
  assign _T_2384 = _T_2378 & auto_in_a_valid; // @[ToAXI4.scala 178:31:boom.system.TestHarness.MegaBoomConfig.fir@20371.4]
  assign _T_2385 = _T_2365 == 1'h0; // @[ToAXI4.scala 178:61:boom.system.TestHarness.MegaBoomConfig.fir@20372.4]
  assign _T_2386 = _T_2385 & _T_2341_ready; // @[ToAXI4.scala 178:69:boom.system.TestHarness.MegaBoomConfig.fir@20373.4]
  assign _T_2387 = _T_2296 ? _T_2386 : 1'h1; // @[ToAXI4.scala 178:51:boom.system.TestHarness.MegaBoomConfig.fir@20374.4]
  assign _T_2388 = _T_2384 & _T_2387; // @[ToAXI4.scala 178:45:boom.system.TestHarness.MegaBoomConfig.fir@20375.4]
  assign _T_2391 = _T_2384 & _T_2296; // @[ToAXI4.scala 180:43:boom.system.TestHarness.MegaBoomConfig.fir@20379.4]
  assign _T_2396 = auto_in_d_ready & auto_out_r_valid; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@20387.4]
  assign _T_2397 = auto_out_r_bits_last == 1'h0; // @[ToAXI4.scala 188:42:boom.system.TestHarness.MegaBoomConfig.fir@20389.6]
  assign _T_2398 = auto_out_r_valid | _T_2395; // @[ToAXI4.scala 190:32:boom.system.TestHarness.MegaBoomConfig.fir@20392.4]
  assign _T_2399 = _T_2398 == 1'h0; // @[ToAXI4.scala 193:36:boom.system.TestHarness.MegaBoomConfig.fir@20394.4]
  assign _T_2401 = _T_2398 ? auto_out_r_valid : auto_out_b_valid; // @[ToAXI4.scala 194:24:boom.system.TestHarness.MegaBoomConfig.fir@20397.4]
  assign _T_2405 = auto_out_r_bits_resp == 2'h3; // @[ToAXI4.scala 201:39:boom.system.TestHarness.MegaBoomConfig.fir@20404.4]
  assign _GEN_516 = _T_2403 ? _T_2405 : _T_2407; // @[Reg.scala 12:19:boom.system.TestHarness.MegaBoomConfig.fir@20406.4]
  assign _T_2409 = auto_out_r_bits_resp != 2'h0; // @[ToAXI4.scala 202:39:boom.system.TestHarness.MegaBoomConfig.fir@20410.4]
  assign _T_2410 = auto_out_b_bits_resp != 2'h0; // @[ToAXI4.scala 203:39:boom.system.TestHarness.MegaBoomConfig.fir@20411.4]
  assign _T_2411 = _T_2409 | _GEN_516; // @[ToAXI4.scala 205:100:boom.system.TestHarness.MegaBoomConfig.fir@20412.4]
  assign _T_2418 = 256'h1 << _GEN_257; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@20437.4]
  assign _T_2420 = _T_2418[0]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20439.4]
  assign _T_2421 = _T_2418[1]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20440.4]
  assign _T_2422 = _T_2418[2]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20441.4]
  assign _T_2423 = _T_2418[3]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20442.4]
  assign _T_2424 = _T_2418[4]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20443.4]
  assign _T_2425 = _T_2418[5]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20444.4]
  assign _T_2426 = _T_2418[6]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20445.4]
  assign _T_2427 = _T_2418[7]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20446.4]
  assign _T_2428 = _T_2418[8]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20447.4]
  assign _T_2429 = _T_2418[9]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20448.4]
  assign _T_2430 = _T_2418[10]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20449.4]
  assign _T_2431 = _T_2418[11]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20450.4]
  assign _T_2432 = _T_2418[12]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20451.4]
  assign _T_2433 = _T_2418[13]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20452.4]
  assign _T_2434 = _T_2418[14]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20453.4]
  assign _T_2435 = _T_2418[15]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20454.4]
  assign _T_2436 = _T_2418[16]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20455.4]
  assign _T_2437 = _T_2418[17]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20456.4]
  assign _T_2438 = _T_2418[18]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20457.4]
  assign _T_2439 = _T_2418[19]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20458.4]
  assign _T_2440 = _T_2418[20]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20459.4]
  assign _T_2441 = _T_2418[21]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20460.4]
  assign _T_2442 = _T_2418[22]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20461.4]
  assign _T_2443 = _T_2418[23]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20462.4]
  assign _T_2444 = _T_2418[24]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20463.4]
  assign _T_2445 = _T_2418[25]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20464.4]
  assign _T_2446 = _T_2418[26]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20465.4]
  assign _T_2447 = _T_2418[27]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20466.4]
  assign _T_2448 = _T_2418[28]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20467.4]
  assign _T_2449 = _T_2418[29]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20468.4]
  assign _T_2450 = _T_2418[30]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20469.4]
  assign _T_2451 = _T_2418[31]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20470.4]
  assign _T_2452 = _T_2418[32]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20471.4]
  assign _T_2453 = _T_2418[33]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20472.4]
  assign _T_2454 = _T_2418[34]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20473.4]
  assign _T_2455 = _T_2418[35]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20474.4]
  assign _T_2456 = _T_2418[36]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20475.4]
  assign _T_2457 = _T_2418[37]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20476.4]
  assign _T_2458 = _T_2418[38]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20477.4]
  assign _T_2459 = _T_2418[39]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20478.4]
  assign _T_2460 = _T_2418[40]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20479.4]
  assign _T_2461 = _T_2418[41]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20480.4]
  assign _T_2462 = _T_2418[42]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20481.4]
  assign _T_2463 = _T_2418[43]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20482.4]
  assign _T_2464 = _T_2418[44]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20483.4]
  assign _T_2465 = _T_2418[45]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20484.4]
  assign _T_2466 = _T_2418[46]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20485.4]
  assign _T_2467 = _T_2418[47]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20486.4]
  assign _T_2468 = _T_2418[48]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20487.4]
  assign _T_2469 = _T_2418[49]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20488.4]
  assign _T_2470 = _T_2418[50]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20489.4]
  assign _T_2471 = _T_2418[51]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20490.4]
  assign _T_2472 = _T_2418[52]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20491.4]
  assign _T_2473 = _T_2418[53]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20492.4]
  assign _T_2474 = _T_2418[54]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20493.4]
  assign _T_2475 = _T_2418[55]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20494.4]
  assign _T_2476 = _T_2418[56]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20495.4]
  assign _T_2477 = _T_2418[57]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20496.4]
  assign _T_2478 = _T_2418[58]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20497.4]
  assign _T_2479 = _T_2418[59]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20498.4]
  assign _T_2480 = _T_2418[60]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20499.4]
  assign _T_2481 = _T_2418[61]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20500.4]
  assign _T_2482 = _T_2418[62]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20501.4]
  assign _T_2483 = _T_2418[63]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20502.4]
  assign _T_2484 = _T_2418[64]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20503.4]
  assign _T_2485 = _T_2418[65]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20504.4]
  assign _T_2486 = _T_2418[66]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20505.4]
  assign _T_2487 = _T_2418[67]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20506.4]
  assign _T_2488 = _T_2418[68]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20507.4]
  assign _T_2489 = _T_2418[69]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20508.4]
  assign _T_2490 = _T_2418[70]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20509.4]
  assign _T_2491 = _T_2418[71]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20510.4]
  assign _T_2492 = _T_2418[72]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20511.4]
  assign _T_2493 = _T_2418[73]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20512.4]
  assign _T_2494 = _T_2418[74]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20513.4]
  assign _T_2495 = _T_2418[75]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20514.4]
  assign _T_2496 = _T_2418[76]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20515.4]
  assign _T_2497 = _T_2418[77]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20516.4]
  assign _T_2498 = _T_2418[78]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20517.4]
  assign _T_2499 = _T_2418[79]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20518.4]
  assign _T_2500 = _T_2418[80]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20519.4]
  assign _T_2501 = _T_2418[81]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20520.4]
  assign _T_2502 = _T_2418[82]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20521.4]
  assign _T_2503 = _T_2418[83]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20522.4]
  assign _T_2504 = _T_2418[84]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20523.4]
  assign _T_2505 = _T_2418[85]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20524.4]
  assign _T_2506 = _T_2418[86]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20525.4]
  assign _T_2507 = _T_2418[87]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20526.4]
  assign _T_2508 = _T_2418[88]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20527.4]
  assign _T_2509 = _T_2418[89]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20528.4]
  assign _T_2510 = _T_2418[90]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20529.4]
  assign _T_2511 = _T_2418[91]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20530.4]
  assign _T_2512 = _T_2418[92]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20531.4]
  assign _T_2513 = _T_2418[93]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20532.4]
  assign _T_2514 = _T_2418[94]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20533.4]
  assign _T_2515 = _T_2418[95]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20534.4]
  assign _T_2516 = _T_2418[96]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20535.4]
  assign _T_2517 = _T_2418[97]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20536.4]
  assign _T_2518 = _T_2418[98]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20537.4]
  assign _T_2519 = _T_2418[99]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20538.4]
  assign _T_2520 = _T_2418[100]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20539.4]
  assign _T_2521 = _T_2418[101]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20540.4]
  assign _T_2522 = _T_2418[102]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20541.4]
  assign _T_2523 = _T_2418[103]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20542.4]
  assign _T_2524 = _T_2418[104]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20543.4]
  assign _T_2525 = _T_2418[105]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20544.4]
  assign _T_2526 = _T_2418[106]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20545.4]
  assign _T_2527 = _T_2418[107]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20546.4]
  assign _T_2528 = _T_2418[108]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20547.4]
  assign _T_2529 = _T_2418[109]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20548.4]
  assign _T_2530 = _T_2418[110]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20549.4]
  assign _T_2531 = _T_2418[111]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20550.4]
  assign _T_2532 = _T_2418[112]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20551.4]
  assign _T_2533 = _T_2418[113]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20552.4]
  assign _T_2534 = _T_2418[114]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20553.4]
  assign _T_2535 = _T_2418[115]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20554.4]
  assign _T_2536 = _T_2418[116]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20555.4]
  assign _T_2537 = _T_2418[117]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20556.4]
  assign _T_2538 = _T_2418[118]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20557.4]
  assign _T_2539 = _T_2418[119]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20558.4]
  assign _T_2540 = _T_2418[120]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20559.4]
  assign _T_2541 = _T_2418[121]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20560.4]
  assign _T_2542 = _T_2418[122]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20561.4]
  assign _T_2543 = _T_2418[123]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20562.4]
  assign _T_2544 = _T_2418[124]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20563.4]
  assign _T_2545 = _T_2418[125]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20564.4]
  assign _T_2546 = _T_2418[126]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20565.4]
  assign _T_2547 = _T_2418[127]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20566.4]
  assign _T_2548 = _T_2418[128]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20567.4]
  assign _T_2549 = _T_2418[129]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20568.4]
  assign _T_2550 = _T_2418[130]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20569.4]
  assign _T_2551 = _T_2418[131]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20570.4]
  assign _T_2552 = _T_2418[132]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20571.4]
  assign _T_2553 = _T_2418[133]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20572.4]
  assign _T_2554 = _T_2418[134]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20573.4]
  assign _T_2555 = _T_2418[135]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20574.4]
  assign _T_2556 = _T_2418[136]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20575.4]
  assign _T_2557 = _T_2418[137]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20576.4]
  assign _T_2558 = _T_2418[138]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20577.4]
  assign _T_2559 = _T_2418[139]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20578.4]
  assign _T_2560 = _T_2418[140]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20579.4]
  assign _T_2561 = _T_2418[141]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20580.4]
  assign _T_2562 = _T_2418[142]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20581.4]
  assign _T_2563 = _T_2418[143]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20582.4]
  assign _T_2564 = _T_2418[144]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20583.4]
  assign _T_2565 = _T_2418[145]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20584.4]
  assign _T_2566 = _T_2418[146]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20585.4]
  assign _T_2567 = _T_2418[147]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20586.4]
  assign _T_2568 = _T_2418[148]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20587.4]
  assign _T_2569 = _T_2418[149]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20588.4]
  assign _T_2570 = _T_2418[150]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20589.4]
  assign _T_2571 = _T_2418[151]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20590.4]
  assign _T_2572 = _T_2418[152]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20591.4]
  assign _T_2573 = _T_2418[153]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20592.4]
  assign _T_2574 = _T_2418[154]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20593.4]
  assign _T_2575 = _T_2418[155]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20594.4]
  assign _T_2576 = _T_2418[156]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20595.4]
  assign _T_2577 = _T_2418[157]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20596.4]
  assign _T_2578 = _T_2418[158]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20597.4]
  assign _T_2579 = _T_2418[159]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20598.4]
  assign _T_2580 = _T_2418[160]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20599.4]
  assign _T_2581 = _T_2418[161]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20600.4]
  assign _T_2582 = _T_2418[162]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20601.4]
  assign _T_2583 = _T_2418[163]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20602.4]
  assign _T_2584 = _T_2418[164]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20603.4]
  assign _T_2585 = _T_2418[165]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20604.4]
  assign _T_2586 = _T_2418[166]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20605.4]
  assign _T_2587 = _T_2418[167]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20606.4]
  assign _T_2588 = _T_2418[168]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20607.4]
  assign _T_2589 = _T_2418[169]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20608.4]
  assign _T_2590 = _T_2418[170]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20609.4]
  assign _T_2591 = _T_2418[171]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20610.4]
  assign _T_2592 = _T_2418[172]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20611.4]
  assign _T_2593 = _T_2418[173]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20612.4]
  assign _T_2594 = _T_2418[174]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20613.4]
  assign _T_2595 = _T_2418[175]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20614.4]
  assign _T_2596 = _T_2418[176]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20615.4]
  assign _T_2597 = _T_2418[177]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20616.4]
  assign _T_2598 = _T_2418[178]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20617.4]
  assign _T_2599 = _T_2418[179]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20618.4]
  assign _T_2600 = _T_2418[180]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20619.4]
  assign _T_2601 = _T_2418[181]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20620.4]
  assign _T_2602 = _T_2418[182]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20621.4]
  assign _T_2603 = _T_2418[183]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20622.4]
  assign _T_2604 = _T_2418[184]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20623.4]
  assign _T_2605 = _T_2418[185]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20624.4]
  assign _T_2606 = _T_2418[186]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20625.4]
  assign _T_2607 = _T_2418[187]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20626.4]
  assign _T_2608 = _T_2418[188]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20627.4]
  assign _T_2609 = _T_2418[189]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20628.4]
  assign _T_2610 = _T_2418[190]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20629.4]
  assign _T_2611 = _T_2418[191]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20630.4]
  assign _T_2612 = _T_2418[192]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20631.4]
  assign _T_2613 = _T_2418[193]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20632.4]
  assign _T_2614 = _T_2418[194]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20633.4]
  assign _T_2615 = _T_2418[195]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20634.4]
  assign _T_2616 = _T_2418[196]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20635.4]
  assign _T_2617 = _T_2418[197]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20636.4]
  assign _T_2618 = _T_2418[198]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20637.4]
  assign _T_2619 = _T_2418[199]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20638.4]
  assign _T_2620 = _T_2418[200]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20639.4]
  assign _T_2621 = _T_2418[201]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20640.4]
  assign _T_2622 = _T_2418[202]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20641.4]
  assign _T_2623 = _T_2418[203]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20642.4]
  assign _T_2624 = _T_2418[204]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20643.4]
  assign _T_2625 = _T_2418[205]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20644.4]
  assign _T_2626 = _T_2418[206]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20645.4]
  assign _T_2627 = _T_2418[207]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20646.4]
  assign _T_2628 = _T_2418[208]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20647.4]
  assign _T_2629 = _T_2418[209]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20648.4]
  assign _T_2630 = _T_2418[210]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20649.4]
  assign _T_2631 = _T_2418[211]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20650.4]
  assign _T_2632 = _T_2418[212]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20651.4]
  assign _T_2633 = _T_2418[213]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20652.4]
  assign _T_2634 = _T_2418[214]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20653.4]
  assign _T_2635 = _T_2418[215]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20654.4]
  assign _T_2636 = _T_2418[216]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20655.4]
  assign _T_2637 = _T_2418[217]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20656.4]
  assign _T_2638 = _T_2418[218]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20657.4]
  assign _T_2639 = _T_2418[219]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20658.4]
  assign _T_2640 = _T_2418[220]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20659.4]
  assign _T_2641 = _T_2418[221]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20660.4]
  assign _T_2642 = _T_2418[222]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20661.4]
  assign _T_2643 = _T_2418[223]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20662.4]
  assign _T_2644 = _T_2418[224]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20663.4]
  assign _T_2645 = _T_2418[225]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20664.4]
  assign _T_2646 = _T_2418[226]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20665.4]
  assign _T_2647 = _T_2418[227]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20666.4]
  assign _T_2648 = _T_2418[228]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20667.4]
  assign _T_2649 = _T_2418[229]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20668.4]
  assign _T_2650 = _T_2418[230]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20669.4]
  assign _T_2651 = _T_2418[231]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20670.4]
  assign _T_2652 = _T_2418[232]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20671.4]
  assign _T_2653 = _T_2418[233]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20672.4]
  assign _T_2654 = _T_2418[234]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20673.4]
  assign _T_2655 = _T_2418[235]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20674.4]
  assign _T_2656 = _T_2418[236]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20675.4]
  assign _T_2657 = _T_2418[237]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20676.4]
  assign _T_2658 = _T_2418[238]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20677.4]
  assign _T_2659 = _T_2418[239]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20678.4]
  assign _T_2660 = _T_2418[240]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20679.4]
  assign _T_2661 = _T_2418[241]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20680.4]
  assign _T_2662 = _T_2418[242]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20681.4]
  assign _T_2663 = _T_2418[243]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20682.4]
  assign _T_2664 = _T_2418[244]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20683.4]
  assign _T_2665 = _T_2418[245]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20684.4]
  assign _T_2666 = _T_2418[246]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20685.4]
  assign _T_2667 = _T_2418[247]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20686.4]
  assign _T_2668 = _T_2418[248]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20687.4]
  assign _T_2669 = _T_2418[249]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20688.4]
  assign _T_2670 = _T_2418[250]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20689.4]
  assign _T_2671 = _T_2418[251]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20690.4]
  assign _T_2672 = _T_2418[252]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20691.4]
  assign _T_2673 = _T_2418[253]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20692.4]
  assign _T_2674 = _T_2418[254]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20693.4]
  assign _T_2675 = _T_2418[255]; // @[ToAXI4.scala 213:58:boom.system.TestHarness.MegaBoomConfig.fir@20694.4]
  assign _T_2676 = _T_2398 ? auto_out_r_bits_id : auto_out_b_bits_id; // @[ToAXI4.scala 214:31:boom.system.TestHarness.MegaBoomConfig.fir@20695.4]
  assign _T_2678 = 256'h1 << _T_2676; // @[OneHot.scala 52:12:boom.system.TestHarness.MegaBoomConfig.fir@20697.4]
  assign _T_2680 = _T_2678[0]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20699.4]
  assign _T_2681 = _T_2678[1]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20700.4]
  assign _T_2682 = _T_2678[2]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20701.4]
  assign _T_2683 = _T_2678[3]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20702.4]
  assign _T_2684 = _T_2678[4]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20703.4]
  assign _T_2685 = _T_2678[5]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20704.4]
  assign _T_2686 = _T_2678[6]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20705.4]
  assign _T_2687 = _T_2678[7]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20706.4]
  assign _T_2688 = _T_2678[8]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20707.4]
  assign _T_2689 = _T_2678[9]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20708.4]
  assign _T_2690 = _T_2678[10]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20709.4]
  assign _T_2691 = _T_2678[11]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20710.4]
  assign _T_2692 = _T_2678[12]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20711.4]
  assign _T_2693 = _T_2678[13]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20712.4]
  assign _T_2694 = _T_2678[14]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20713.4]
  assign _T_2695 = _T_2678[15]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20714.4]
  assign _T_2696 = _T_2678[16]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20715.4]
  assign _T_2697 = _T_2678[17]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20716.4]
  assign _T_2698 = _T_2678[18]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20717.4]
  assign _T_2699 = _T_2678[19]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20718.4]
  assign _T_2700 = _T_2678[20]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20719.4]
  assign _T_2701 = _T_2678[21]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20720.4]
  assign _T_2702 = _T_2678[22]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20721.4]
  assign _T_2703 = _T_2678[23]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20722.4]
  assign _T_2704 = _T_2678[24]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20723.4]
  assign _T_2705 = _T_2678[25]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20724.4]
  assign _T_2706 = _T_2678[26]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20725.4]
  assign _T_2707 = _T_2678[27]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20726.4]
  assign _T_2708 = _T_2678[28]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20727.4]
  assign _T_2709 = _T_2678[29]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20728.4]
  assign _T_2710 = _T_2678[30]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20729.4]
  assign _T_2711 = _T_2678[31]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20730.4]
  assign _T_2712 = _T_2678[32]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20731.4]
  assign _T_2713 = _T_2678[33]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20732.4]
  assign _T_2714 = _T_2678[34]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20733.4]
  assign _T_2715 = _T_2678[35]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20734.4]
  assign _T_2716 = _T_2678[36]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20735.4]
  assign _T_2717 = _T_2678[37]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20736.4]
  assign _T_2718 = _T_2678[38]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20737.4]
  assign _T_2719 = _T_2678[39]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20738.4]
  assign _T_2720 = _T_2678[40]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20739.4]
  assign _T_2721 = _T_2678[41]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20740.4]
  assign _T_2722 = _T_2678[42]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20741.4]
  assign _T_2723 = _T_2678[43]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20742.4]
  assign _T_2724 = _T_2678[44]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20743.4]
  assign _T_2725 = _T_2678[45]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20744.4]
  assign _T_2726 = _T_2678[46]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20745.4]
  assign _T_2727 = _T_2678[47]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20746.4]
  assign _T_2728 = _T_2678[48]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20747.4]
  assign _T_2729 = _T_2678[49]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20748.4]
  assign _T_2730 = _T_2678[50]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20749.4]
  assign _T_2731 = _T_2678[51]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20750.4]
  assign _T_2732 = _T_2678[52]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20751.4]
  assign _T_2733 = _T_2678[53]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20752.4]
  assign _T_2734 = _T_2678[54]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20753.4]
  assign _T_2735 = _T_2678[55]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20754.4]
  assign _T_2736 = _T_2678[56]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20755.4]
  assign _T_2737 = _T_2678[57]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20756.4]
  assign _T_2738 = _T_2678[58]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20757.4]
  assign _T_2739 = _T_2678[59]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20758.4]
  assign _T_2740 = _T_2678[60]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20759.4]
  assign _T_2741 = _T_2678[61]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20760.4]
  assign _T_2742 = _T_2678[62]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20761.4]
  assign _T_2743 = _T_2678[63]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20762.4]
  assign _T_2744 = _T_2678[64]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20763.4]
  assign _T_2745 = _T_2678[65]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20764.4]
  assign _T_2746 = _T_2678[66]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20765.4]
  assign _T_2747 = _T_2678[67]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20766.4]
  assign _T_2748 = _T_2678[68]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20767.4]
  assign _T_2749 = _T_2678[69]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20768.4]
  assign _T_2750 = _T_2678[70]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20769.4]
  assign _T_2751 = _T_2678[71]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20770.4]
  assign _T_2752 = _T_2678[72]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20771.4]
  assign _T_2753 = _T_2678[73]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20772.4]
  assign _T_2754 = _T_2678[74]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20773.4]
  assign _T_2755 = _T_2678[75]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20774.4]
  assign _T_2756 = _T_2678[76]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20775.4]
  assign _T_2757 = _T_2678[77]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20776.4]
  assign _T_2758 = _T_2678[78]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20777.4]
  assign _T_2759 = _T_2678[79]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20778.4]
  assign _T_2760 = _T_2678[80]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20779.4]
  assign _T_2761 = _T_2678[81]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20780.4]
  assign _T_2762 = _T_2678[82]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20781.4]
  assign _T_2763 = _T_2678[83]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20782.4]
  assign _T_2764 = _T_2678[84]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20783.4]
  assign _T_2765 = _T_2678[85]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20784.4]
  assign _T_2766 = _T_2678[86]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20785.4]
  assign _T_2767 = _T_2678[87]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20786.4]
  assign _T_2768 = _T_2678[88]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20787.4]
  assign _T_2769 = _T_2678[89]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20788.4]
  assign _T_2770 = _T_2678[90]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20789.4]
  assign _T_2771 = _T_2678[91]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20790.4]
  assign _T_2772 = _T_2678[92]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20791.4]
  assign _T_2773 = _T_2678[93]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20792.4]
  assign _T_2774 = _T_2678[94]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20793.4]
  assign _T_2775 = _T_2678[95]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20794.4]
  assign _T_2776 = _T_2678[96]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20795.4]
  assign _T_2777 = _T_2678[97]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20796.4]
  assign _T_2778 = _T_2678[98]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20797.4]
  assign _T_2779 = _T_2678[99]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20798.4]
  assign _T_2780 = _T_2678[100]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20799.4]
  assign _T_2781 = _T_2678[101]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20800.4]
  assign _T_2782 = _T_2678[102]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20801.4]
  assign _T_2783 = _T_2678[103]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20802.4]
  assign _T_2784 = _T_2678[104]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20803.4]
  assign _T_2785 = _T_2678[105]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20804.4]
  assign _T_2786 = _T_2678[106]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20805.4]
  assign _T_2787 = _T_2678[107]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20806.4]
  assign _T_2788 = _T_2678[108]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20807.4]
  assign _T_2789 = _T_2678[109]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20808.4]
  assign _T_2790 = _T_2678[110]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20809.4]
  assign _T_2791 = _T_2678[111]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20810.4]
  assign _T_2792 = _T_2678[112]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20811.4]
  assign _T_2793 = _T_2678[113]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20812.4]
  assign _T_2794 = _T_2678[114]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20813.4]
  assign _T_2795 = _T_2678[115]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20814.4]
  assign _T_2796 = _T_2678[116]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20815.4]
  assign _T_2797 = _T_2678[117]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20816.4]
  assign _T_2798 = _T_2678[118]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20817.4]
  assign _T_2799 = _T_2678[119]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20818.4]
  assign _T_2800 = _T_2678[120]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20819.4]
  assign _T_2801 = _T_2678[121]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20820.4]
  assign _T_2802 = _T_2678[122]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20821.4]
  assign _T_2803 = _T_2678[123]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20822.4]
  assign _T_2804 = _T_2678[124]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20823.4]
  assign _T_2805 = _T_2678[125]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20824.4]
  assign _T_2806 = _T_2678[126]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20825.4]
  assign _T_2807 = _T_2678[127]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20826.4]
  assign _T_2808 = _T_2678[128]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20827.4]
  assign _T_2809 = _T_2678[129]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20828.4]
  assign _T_2810 = _T_2678[130]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20829.4]
  assign _T_2811 = _T_2678[131]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20830.4]
  assign _T_2812 = _T_2678[132]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20831.4]
  assign _T_2813 = _T_2678[133]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20832.4]
  assign _T_2814 = _T_2678[134]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20833.4]
  assign _T_2815 = _T_2678[135]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20834.4]
  assign _T_2816 = _T_2678[136]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20835.4]
  assign _T_2817 = _T_2678[137]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20836.4]
  assign _T_2818 = _T_2678[138]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20837.4]
  assign _T_2819 = _T_2678[139]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20838.4]
  assign _T_2820 = _T_2678[140]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20839.4]
  assign _T_2821 = _T_2678[141]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20840.4]
  assign _T_2822 = _T_2678[142]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20841.4]
  assign _T_2823 = _T_2678[143]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20842.4]
  assign _T_2824 = _T_2678[144]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20843.4]
  assign _T_2825 = _T_2678[145]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20844.4]
  assign _T_2826 = _T_2678[146]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20845.4]
  assign _T_2827 = _T_2678[147]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20846.4]
  assign _T_2828 = _T_2678[148]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20847.4]
  assign _T_2829 = _T_2678[149]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20848.4]
  assign _T_2830 = _T_2678[150]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20849.4]
  assign _T_2831 = _T_2678[151]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20850.4]
  assign _T_2832 = _T_2678[152]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20851.4]
  assign _T_2833 = _T_2678[153]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20852.4]
  assign _T_2834 = _T_2678[154]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20853.4]
  assign _T_2835 = _T_2678[155]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20854.4]
  assign _T_2836 = _T_2678[156]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20855.4]
  assign _T_2837 = _T_2678[157]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20856.4]
  assign _T_2838 = _T_2678[158]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20857.4]
  assign _T_2839 = _T_2678[159]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20858.4]
  assign _T_2840 = _T_2678[160]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20859.4]
  assign _T_2841 = _T_2678[161]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20860.4]
  assign _T_2842 = _T_2678[162]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20861.4]
  assign _T_2843 = _T_2678[163]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20862.4]
  assign _T_2844 = _T_2678[164]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20863.4]
  assign _T_2845 = _T_2678[165]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20864.4]
  assign _T_2846 = _T_2678[166]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20865.4]
  assign _T_2847 = _T_2678[167]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20866.4]
  assign _T_2848 = _T_2678[168]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20867.4]
  assign _T_2849 = _T_2678[169]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20868.4]
  assign _T_2850 = _T_2678[170]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20869.4]
  assign _T_2851 = _T_2678[171]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20870.4]
  assign _T_2852 = _T_2678[172]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20871.4]
  assign _T_2853 = _T_2678[173]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20872.4]
  assign _T_2854 = _T_2678[174]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20873.4]
  assign _T_2855 = _T_2678[175]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20874.4]
  assign _T_2856 = _T_2678[176]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20875.4]
  assign _T_2857 = _T_2678[177]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20876.4]
  assign _T_2858 = _T_2678[178]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20877.4]
  assign _T_2859 = _T_2678[179]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20878.4]
  assign _T_2860 = _T_2678[180]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20879.4]
  assign _T_2861 = _T_2678[181]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20880.4]
  assign _T_2862 = _T_2678[182]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20881.4]
  assign _T_2863 = _T_2678[183]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20882.4]
  assign _T_2864 = _T_2678[184]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20883.4]
  assign _T_2865 = _T_2678[185]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20884.4]
  assign _T_2866 = _T_2678[186]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20885.4]
  assign _T_2867 = _T_2678[187]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20886.4]
  assign _T_2868 = _T_2678[188]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20887.4]
  assign _T_2869 = _T_2678[189]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20888.4]
  assign _T_2870 = _T_2678[190]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20889.4]
  assign _T_2871 = _T_2678[191]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20890.4]
  assign _T_2872 = _T_2678[192]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20891.4]
  assign _T_2873 = _T_2678[193]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20892.4]
  assign _T_2874 = _T_2678[194]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20893.4]
  assign _T_2875 = _T_2678[195]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20894.4]
  assign _T_2876 = _T_2678[196]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20895.4]
  assign _T_2877 = _T_2678[197]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20896.4]
  assign _T_2878 = _T_2678[198]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20897.4]
  assign _T_2879 = _T_2678[199]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20898.4]
  assign _T_2880 = _T_2678[200]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20899.4]
  assign _T_2881 = _T_2678[201]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20900.4]
  assign _T_2882 = _T_2678[202]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20901.4]
  assign _T_2883 = _T_2678[203]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20902.4]
  assign _T_2884 = _T_2678[204]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20903.4]
  assign _T_2885 = _T_2678[205]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20904.4]
  assign _T_2886 = _T_2678[206]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20905.4]
  assign _T_2887 = _T_2678[207]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20906.4]
  assign _T_2888 = _T_2678[208]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20907.4]
  assign _T_2889 = _T_2678[209]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20908.4]
  assign _T_2890 = _T_2678[210]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20909.4]
  assign _T_2891 = _T_2678[211]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20910.4]
  assign _T_2892 = _T_2678[212]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20911.4]
  assign _T_2893 = _T_2678[213]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20912.4]
  assign _T_2894 = _T_2678[214]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20913.4]
  assign _T_2895 = _T_2678[215]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20914.4]
  assign _T_2896 = _T_2678[216]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20915.4]
  assign _T_2897 = _T_2678[217]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20916.4]
  assign _T_2898 = _T_2678[218]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20917.4]
  assign _T_2899 = _T_2678[219]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20918.4]
  assign _T_2900 = _T_2678[220]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20919.4]
  assign _T_2901 = _T_2678[221]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20920.4]
  assign _T_2902 = _T_2678[222]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20921.4]
  assign _T_2903 = _T_2678[223]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20922.4]
  assign _T_2904 = _T_2678[224]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20923.4]
  assign _T_2905 = _T_2678[225]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20924.4]
  assign _T_2906 = _T_2678[226]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20925.4]
  assign _T_2907 = _T_2678[227]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20926.4]
  assign _T_2908 = _T_2678[228]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20927.4]
  assign _T_2909 = _T_2678[229]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20928.4]
  assign _T_2910 = _T_2678[230]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20929.4]
  assign _T_2911 = _T_2678[231]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20930.4]
  assign _T_2912 = _T_2678[232]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20931.4]
  assign _T_2913 = _T_2678[233]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20932.4]
  assign _T_2914 = _T_2678[234]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20933.4]
  assign _T_2915 = _T_2678[235]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20934.4]
  assign _T_2916 = _T_2678[236]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20935.4]
  assign _T_2917 = _T_2678[237]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20936.4]
  assign _T_2918 = _T_2678[238]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20937.4]
  assign _T_2919 = _T_2678[239]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20938.4]
  assign _T_2920 = _T_2678[240]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20939.4]
  assign _T_2921 = _T_2678[241]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20940.4]
  assign _T_2922 = _T_2678[242]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20941.4]
  assign _T_2923 = _T_2678[243]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20942.4]
  assign _T_2924 = _T_2678[244]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20943.4]
  assign _T_2925 = _T_2678[245]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20944.4]
  assign _T_2926 = _T_2678[246]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20945.4]
  assign _T_2927 = _T_2678[247]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20946.4]
  assign _T_2928 = _T_2678[248]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20947.4]
  assign _T_2929 = _T_2678[249]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20948.4]
  assign _T_2930 = _T_2678[250]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20949.4]
  assign _T_2931 = _T_2678[251]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20950.4]
  assign _T_2932 = _T_2678[252]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20951.4]
  assign _T_2933 = _T_2678[253]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20952.4]
  assign _T_2934 = _T_2678[254]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20953.4]
  assign _T_2935 = _T_2678[255]; // @[ToAXI4.scala 214:93:boom.system.TestHarness.MegaBoomConfig.fir@20954.4]
  assign _T_2936 = _T_2398 ? auto_out_r_bits_last : 1'h1; // @[ToAXI4.scala 215:23:boom.system.TestHarness.MegaBoomConfig.fir@20955.4]
  assign _T_2942 = _T_2338_ready & _T_2388; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@20959.4]
  assign _T_2943 = _T_2420 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@20960.4]
  assign _T_2944 = _T_2680 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@20961.4]
  assign _T_2945 = auto_in_d_ready & _T_2401; // @[Decoupled.scala 37:37:boom.system.TestHarness.MegaBoomConfig.fir@20962.4]
  assign _T_2946 = _T_2944 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@20963.4]
  assign _T_2948 = _T_2938 + _T_2943; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@20965.4]
  assign _T_2949 = _T_2948 - _T_2946; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@20966.4]
  assign _T_2950 = $unsigned(_T_2949); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@20967.4]
  assign _T_2951 = _T_2950[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@20968.4]
  assign _T_2952 = _T_2946 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@20970.4]
  assign _T_2954 = _T_2952 | _T_2938; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@20972.4]
  assign _T_2956 = _T_2954 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@20974.4]
  assign _T_2957 = _T_2956 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@20975.4]
  assign _T_2958 = _T_2943 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@20980.4]
  assign _T_2959 = _T_2938 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@20981.4]
  assign _T_2960 = _T_2958 | _T_2959; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@20982.4]
  assign _T_2962 = _T_2960 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@20984.4]
  assign _T_2963 = _T_2962 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@20985.4]
  assign _T_2974 = _T_2421 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21002.4]
  assign _T_2975 = _T_2681 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21003.4]
  assign _T_2977 = _T_2975 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21005.4]
  assign _T_2979 = _T_2969 + _T_2974; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21007.4]
  assign _T_2980 = _T_2979 - _T_2977; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21008.4]
  assign _T_2981 = $unsigned(_T_2980); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21009.4]
  assign _T_2982 = _T_2981[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21010.4]
  assign _T_2983 = _T_2977 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21012.4]
  assign _T_2985 = _T_2983 | _T_2969; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21014.4]
  assign _T_2987 = _T_2985 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21016.4]
  assign _T_2988 = _T_2987 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21017.4]
  assign _T_2989 = _T_2974 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21022.4]
  assign _T_2990 = _T_2969 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21023.4]
  assign _T_2991 = _T_2989 | _T_2990; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21024.4]
  assign _T_2993 = _T_2991 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21026.4]
  assign _T_2994 = _T_2993 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21027.4]
  assign _T_3005 = _T_2422 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21044.4]
  assign _T_3006 = _T_2682 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21045.4]
  assign _T_3008 = _T_3006 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21047.4]
  assign _T_3010 = _T_3000 + _T_3005; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21049.4]
  assign _T_3011 = _T_3010 - _T_3008; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21050.4]
  assign _T_3012 = $unsigned(_T_3011); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21051.4]
  assign _T_3013 = _T_3012[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21052.4]
  assign _T_3014 = _T_3008 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21054.4]
  assign _T_3016 = _T_3014 | _T_3000; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21056.4]
  assign _T_3018 = _T_3016 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21058.4]
  assign _T_3019 = _T_3018 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21059.4]
  assign _T_3020 = _T_3005 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21064.4]
  assign _T_3021 = _T_3000 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21065.4]
  assign _T_3022 = _T_3020 | _T_3021; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21066.4]
  assign _T_3024 = _T_3022 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21068.4]
  assign _T_3025 = _T_3024 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21069.4]
  assign _T_3036 = _T_2423 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21086.4]
  assign _T_3037 = _T_2683 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21087.4]
  assign _T_3039 = _T_3037 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21089.4]
  assign _T_3041 = _T_3031 + _T_3036; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21091.4]
  assign _T_3042 = _T_3041 - _T_3039; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21092.4]
  assign _T_3043 = $unsigned(_T_3042); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21093.4]
  assign _T_3044 = _T_3043[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21094.4]
  assign _T_3045 = _T_3039 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21096.4]
  assign _T_3047 = _T_3045 | _T_3031; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21098.4]
  assign _T_3049 = _T_3047 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21100.4]
  assign _T_3050 = _T_3049 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21101.4]
  assign _T_3051 = _T_3036 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21106.4]
  assign _T_3052 = _T_3031 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21107.4]
  assign _T_3053 = _T_3051 | _T_3052; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21108.4]
  assign _T_3055 = _T_3053 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21110.4]
  assign _T_3056 = _T_3055 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21111.4]
  assign _T_3067 = _T_2424 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21128.4]
  assign _T_3068 = _T_2684 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21129.4]
  assign _T_3070 = _T_3068 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21131.4]
  assign _T_3072 = _T_3062 + _T_3067; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21133.4]
  assign _T_3073 = _T_3072 - _T_3070; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21134.4]
  assign _T_3074 = $unsigned(_T_3073); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21135.4]
  assign _T_3075 = _T_3074[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21136.4]
  assign _T_3076 = _T_3070 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21138.4]
  assign _T_3078 = _T_3076 | _T_3062; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21140.4]
  assign _T_3080 = _T_3078 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21142.4]
  assign _T_3081 = _T_3080 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21143.4]
  assign _T_3082 = _T_3067 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21148.4]
  assign _T_3083 = _T_3062 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21149.4]
  assign _T_3084 = _T_3082 | _T_3083; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21150.4]
  assign _T_3086 = _T_3084 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21152.4]
  assign _T_3087 = _T_3086 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21153.4]
  assign _T_3098 = _T_2425 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21170.4]
  assign _T_3099 = _T_2685 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21171.4]
  assign _T_3101 = _T_3099 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21173.4]
  assign _T_3103 = _T_3093 + _T_3098; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21175.4]
  assign _T_3104 = _T_3103 - _T_3101; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21176.4]
  assign _T_3105 = $unsigned(_T_3104); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21177.4]
  assign _T_3106 = _T_3105[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21178.4]
  assign _T_3107 = _T_3101 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21180.4]
  assign _T_3109 = _T_3107 | _T_3093; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21182.4]
  assign _T_3111 = _T_3109 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21184.4]
  assign _T_3112 = _T_3111 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21185.4]
  assign _T_3113 = _T_3098 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21190.4]
  assign _T_3114 = _T_3093 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21191.4]
  assign _T_3115 = _T_3113 | _T_3114; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21192.4]
  assign _T_3117 = _T_3115 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21194.4]
  assign _T_3118 = _T_3117 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21195.4]
  assign _T_3129 = _T_2426 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21212.4]
  assign _T_3130 = _T_2686 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21213.4]
  assign _T_3132 = _T_3130 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21215.4]
  assign _T_3134 = _T_3124 + _T_3129; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21217.4]
  assign _T_3135 = _T_3134 - _T_3132; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21218.4]
  assign _T_3136 = $unsigned(_T_3135); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21219.4]
  assign _T_3137 = _T_3136[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21220.4]
  assign _T_3138 = _T_3132 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21222.4]
  assign _T_3140 = _T_3138 | _T_3124; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21224.4]
  assign _T_3142 = _T_3140 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21226.4]
  assign _T_3143 = _T_3142 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21227.4]
  assign _T_3144 = _T_3129 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21232.4]
  assign _T_3145 = _T_3124 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21233.4]
  assign _T_3146 = _T_3144 | _T_3145; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21234.4]
  assign _T_3148 = _T_3146 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21236.4]
  assign _T_3149 = _T_3148 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21237.4]
  assign _T_3160 = _T_2427 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21254.4]
  assign _T_3161 = _T_2687 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21255.4]
  assign _T_3163 = _T_3161 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21257.4]
  assign _T_3165 = _T_3155 + _T_3160; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21259.4]
  assign _T_3166 = _T_3165 - _T_3163; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21260.4]
  assign _T_3167 = $unsigned(_T_3166); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21261.4]
  assign _T_3168 = _T_3167[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21262.4]
  assign _T_3169 = _T_3163 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21264.4]
  assign _T_3171 = _T_3169 | _T_3155; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21266.4]
  assign _T_3173 = _T_3171 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21268.4]
  assign _T_3174 = _T_3173 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21269.4]
  assign _T_3175 = _T_3160 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21274.4]
  assign _T_3176 = _T_3155 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21275.4]
  assign _T_3177 = _T_3175 | _T_3176; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21276.4]
  assign _T_3179 = _T_3177 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21278.4]
  assign _T_3180 = _T_3179 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21279.4]
  assign _T_3191 = _T_2428 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21296.4]
  assign _T_3192 = _T_2688 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21297.4]
  assign _T_3194 = _T_3192 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21299.4]
  assign _T_3196 = _T_3186 + _T_3191; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21301.4]
  assign _T_3197 = _T_3196 - _T_3194; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21302.4]
  assign _T_3198 = $unsigned(_T_3197); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21303.4]
  assign _T_3199 = _T_3198[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21304.4]
  assign _T_3200 = _T_3194 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21306.4]
  assign _T_3202 = _T_3200 | _T_3186; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21308.4]
  assign _T_3204 = _T_3202 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21310.4]
  assign _T_3205 = _T_3204 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21311.4]
  assign _T_3206 = _T_3191 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21316.4]
  assign _T_3207 = _T_3186 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21317.4]
  assign _T_3208 = _T_3206 | _T_3207; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21318.4]
  assign _T_3210 = _T_3208 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21320.4]
  assign _T_3211 = _T_3210 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21321.4]
  assign _T_3222 = _T_2429 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21338.4]
  assign _T_3223 = _T_2689 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21339.4]
  assign _T_3225 = _T_3223 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21341.4]
  assign _T_3227 = _T_3217 + _T_3222; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21343.4]
  assign _T_3228 = _T_3227 - _T_3225; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21344.4]
  assign _T_3229 = $unsigned(_T_3228); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21345.4]
  assign _T_3230 = _T_3229[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21346.4]
  assign _T_3231 = _T_3225 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21348.4]
  assign _T_3233 = _T_3231 | _T_3217; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21350.4]
  assign _T_3235 = _T_3233 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21352.4]
  assign _T_3236 = _T_3235 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21353.4]
  assign _T_3237 = _T_3222 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21358.4]
  assign _T_3238 = _T_3217 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21359.4]
  assign _T_3239 = _T_3237 | _T_3238; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21360.4]
  assign _T_3241 = _T_3239 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21362.4]
  assign _T_3242 = _T_3241 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21363.4]
  assign _T_3253 = _T_2430 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21380.4]
  assign _T_3254 = _T_2690 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21381.4]
  assign _T_3256 = _T_3254 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21383.4]
  assign _T_3258 = _T_3248 + _T_3253; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21385.4]
  assign _T_3259 = _T_3258 - _T_3256; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21386.4]
  assign _T_3260 = $unsigned(_T_3259); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21387.4]
  assign _T_3261 = _T_3260[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21388.4]
  assign _T_3262 = _T_3256 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21390.4]
  assign _T_3264 = _T_3262 | _T_3248; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21392.4]
  assign _T_3266 = _T_3264 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21394.4]
  assign _T_3267 = _T_3266 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21395.4]
  assign _T_3268 = _T_3253 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21400.4]
  assign _T_3269 = _T_3248 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21401.4]
  assign _T_3270 = _T_3268 | _T_3269; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21402.4]
  assign _T_3272 = _T_3270 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21404.4]
  assign _T_3273 = _T_3272 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21405.4]
  assign _T_3284 = _T_2431 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21422.4]
  assign _T_3285 = _T_2691 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21423.4]
  assign _T_3287 = _T_3285 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21425.4]
  assign _T_3289 = _T_3279 + _T_3284; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21427.4]
  assign _T_3290 = _T_3289 - _T_3287; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21428.4]
  assign _T_3291 = $unsigned(_T_3290); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21429.4]
  assign _T_3292 = _T_3291[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21430.4]
  assign _T_3293 = _T_3287 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21432.4]
  assign _T_3295 = _T_3293 | _T_3279; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21434.4]
  assign _T_3297 = _T_3295 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21436.4]
  assign _T_3298 = _T_3297 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21437.4]
  assign _T_3299 = _T_3284 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21442.4]
  assign _T_3300 = _T_3279 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21443.4]
  assign _T_3301 = _T_3299 | _T_3300; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21444.4]
  assign _T_3303 = _T_3301 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21446.4]
  assign _T_3304 = _T_3303 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21447.4]
  assign _T_3315 = _T_2432 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21464.4]
  assign _T_3316 = _T_2692 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21465.4]
  assign _T_3318 = _T_3316 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21467.4]
  assign _T_3320 = _T_3310 + _T_3315; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21469.4]
  assign _T_3321 = _T_3320 - _T_3318; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21470.4]
  assign _T_3322 = $unsigned(_T_3321); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21471.4]
  assign _T_3323 = _T_3322[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21472.4]
  assign _T_3324 = _T_3318 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21474.4]
  assign _T_3326 = _T_3324 | _T_3310; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21476.4]
  assign _T_3328 = _T_3326 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21478.4]
  assign _T_3329 = _T_3328 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21479.4]
  assign _T_3330 = _T_3315 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21484.4]
  assign _T_3331 = _T_3310 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21485.4]
  assign _T_3332 = _T_3330 | _T_3331; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21486.4]
  assign _T_3334 = _T_3332 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21488.4]
  assign _T_3335 = _T_3334 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21489.4]
  assign _T_3346 = _T_2433 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21506.4]
  assign _T_3347 = _T_2693 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21507.4]
  assign _T_3349 = _T_3347 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21509.4]
  assign _T_3351 = _T_3341 + _T_3346; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21511.4]
  assign _T_3352 = _T_3351 - _T_3349; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21512.4]
  assign _T_3353 = $unsigned(_T_3352); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21513.4]
  assign _T_3354 = _T_3353[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21514.4]
  assign _T_3355 = _T_3349 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21516.4]
  assign _T_3357 = _T_3355 | _T_3341; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21518.4]
  assign _T_3359 = _T_3357 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21520.4]
  assign _T_3360 = _T_3359 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21521.4]
  assign _T_3361 = _T_3346 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21526.4]
  assign _T_3362 = _T_3341 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21527.4]
  assign _T_3363 = _T_3361 | _T_3362; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21528.4]
  assign _T_3365 = _T_3363 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21530.4]
  assign _T_3366 = _T_3365 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21531.4]
  assign _T_3377 = _T_2434 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21548.4]
  assign _T_3378 = _T_2694 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21549.4]
  assign _T_3380 = _T_3378 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21551.4]
  assign _T_3382 = _T_3372 + _T_3377; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21553.4]
  assign _T_3383 = _T_3382 - _T_3380; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21554.4]
  assign _T_3384 = $unsigned(_T_3383); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21555.4]
  assign _T_3385 = _T_3384[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21556.4]
  assign _T_3386 = _T_3380 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21558.4]
  assign _T_3388 = _T_3386 | _T_3372; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21560.4]
  assign _T_3390 = _T_3388 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21562.4]
  assign _T_3391 = _T_3390 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21563.4]
  assign _T_3392 = _T_3377 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21568.4]
  assign _T_3393 = _T_3372 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21569.4]
  assign _T_3394 = _T_3392 | _T_3393; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21570.4]
  assign _T_3396 = _T_3394 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21572.4]
  assign _T_3397 = _T_3396 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21573.4]
  assign _T_3408 = _T_2435 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21590.4]
  assign _T_3409 = _T_2695 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21591.4]
  assign _T_3411 = _T_3409 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21593.4]
  assign _T_3413 = _T_3403 + _T_3408; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21595.4]
  assign _T_3414 = _T_3413 - _T_3411; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21596.4]
  assign _T_3415 = $unsigned(_T_3414); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21597.4]
  assign _T_3416 = _T_3415[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21598.4]
  assign _T_3417 = _T_3411 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21600.4]
  assign _T_3419 = _T_3417 | _T_3403; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21602.4]
  assign _T_3421 = _T_3419 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21604.4]
  assign _T_3422 = _T_3421 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21605.4]
  assign _T_3423 = _T_3408 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21610.4]
  assign _T_3424 = _T_3403 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21611.4]
  assign _T_3425 = _T_3423 | _T_3424; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21612.4]
  assign _T_3427 = _T_3425 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21614.4]
  assign _T_3428 = _T_3427 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21615.4]
  assign _T_3439 = _T_2436 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21632.4]
  assign _T_3440 = _T_2696 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21633.4]
  assign _T_3442 = _T_3440 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21635.4]
  assign _T_3444 = _T_3434 + _T_3439; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21637.4]
  assign _T_3445 = _T_3444 - _T_3442; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21638.4]
  assign _T_3446 = $unsigned(_T_3445); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21639.4]
  assign _T_3447 = _T_3446[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21640.4]
  assign _T_3448 = _T_3442 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21642.4]
  assign _T_3450 = _T_3448 | _T_3434; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21644.4]
  assign _T_3452 = _T_3450 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21646.4]
  assign _T_3453 = _T_3452 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21647.4]
  assign _T_3454 = _T_3439 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21652.4]
  assign _T_3455 = _T_3434 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21653.4]
  assign _T_3456 = _T_3454 | _T_3455; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21654.4]
  assign _T_3458 = _T_3456 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21656.4]
  assign _T_3459 = _T_3458 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21657.4]
  assign _T_3470 = _T_2437 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21674.4]
  assign _T_3471 = _T_2697 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21675.4]
  assign _T_3473 = _T_3471 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21677.4]
  assign _T_3475 = _T_3465 + _T_3470; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21679.4]
  assign _T_3476 = _T_3475 - _T_3473; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21680.4]
  assign _T_3477 = $unsigned(_T_3476); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21681.4]
  assign _T_3478 = _T_3477[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21682.4]
  assign _T_3479 = _T_3473 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21684.4]
  assign _T_3481 = _T_3479 | _T_3465; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21686.4]
  assign _T_3483 = _T_3481 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21688.4]
  assign _T_3484 = _T_3483 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21689.4]
  assign _T_3485 = _T_3470 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21694.4]
  assign _T_3486 = _T_3465 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21695.4]
  assign _T_3487 = _T_3485 | _T_3486; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21696.4]
  assign _T_3489 = _T_3487 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21698.4]
  assign _T_3490 = _T_3489 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21699.4]
  assign _T_3501 = _T_2438 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21716.4]
  assign _T_3502 = _T_2698 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21717.4]
  assign _T_3504 = _T_3502 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21719.4]
  assign _T_3506 = _T_3496 + _T_3501; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21721.4]
  assign _T_3507 = _T_3506 - _T_3504; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21722.4]
  assign _T_3508 = $unsigned(_T_3507); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21723.4]
  assign _T_3509 = _T_3508[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21724.4]
  assign _T_3510 = _T_3504 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21726.4]
  assign _T_3512 = _T_3510 | _T_3496; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21728.4]
  assign _T_3514 = _T_3512 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21730.4]
  assign _T_3515 = _T_3514 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21731.4]
  assign _T_3516 = _T_3501 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21736.4]
  assign _T_3517 = _T_3496 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21737.4]
  assign _T_3518 = _T_3516 | _T_3517; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21738.4]
  assign _T_3520 = _T_3518 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21740.4]
  assign _T_3521 = _T_3520 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21741.4]
  assign _T_3532 = _T_2439 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21758.4]
  assign _T_3533 = _T_2699 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21759.4]
  assign _T_3535 = _T_3533 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21761.4]
  assign _T_3537 = _T_3527 + _T_3532; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21763.4]
  assign _T_3538 = _T_3537 - _T_3535; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21764.4]
  assign _T_3539 = $unsigned(_T_3538); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21765.4]
  assign _T_3540 = _T_3539[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21766.4]
  assign _T_3541 = _T_3535 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21768.4]
  assign _T_3543 = _T_3541 | _T_3527; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21770.4]
  assign _T_3545 = _T_3543 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21772.4]
  assign _T_3546 = _T_3545 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21773.4]
  assign _T_3547 = _T_3532 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21778.4]
  assign _T_3548 = _T_3527 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21779.4]
  assign _T_3549 = _T_3547 | _T_3548; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21780.4]
  assign _T_3551 = _T_3549 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21782.4]
  assign _T_3552 = _T_3551 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21783.4]
  assign _T_3563 = _T_2440 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21800.4]
  assign _T_3564 = _T_2700 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21801.4]
  assign _T_3566 = _T_3564 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21803.4]
  assign _T_3568 = _T_3558 + _T_3563; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21805.4]
  assign _T_3569 = _T_3568 - _T_3566; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21806.4]
  assign _T_3570 = $unsigned(_T_3569); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21807.4]
  assign _T_3571 = _T_3570[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21808.4]
  assign _T_3572 = _T_3566 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21810.4]
  assign _T_3574 = _T_3572 | _T_3558; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21812.4]
  assign _T_3576 = _T_3574 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21814.4]
  assign _T_3577 = _T_3576 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21815.4]
  assign _T_3578 = _T_3563 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21820.4]
  assign _T_3579 = _T_3558 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21821.4]
  assign _T_3580 = _T_3578 | _T_3579; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21822.4]
  assign _T_3582 = _T_3580 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21824.4]
  assign _T_3583 = _T_3582 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21825.4]
  assign _T_3594 = _T_2441 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21842.4]
  assign _T_3595 = _T_2701 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21843.4]
  assign _T_3597 = _T_3595 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21845.4]
  assign _T_3599 = _T_3589 + _T_3594; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21847.4]
  assign _T_3600 = _T_3599 - _T_3597; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21848.4]
  assign _T_3601 = $unsigned(_T_3600); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21849.4]
  assign _T_3602 = _T_3601[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21850.4]
  assign _T_3603 = _T_3597 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21852.4]
  assign _T_3605 = _T_3603 | _T_3589; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21854.4]
  assign _T_3607 = _T_3605 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21856.4]
  assign _T_3608 = _T_3607 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21857.4]
  assign _T_3609 = _T_3594 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21862.4]
  assign _T_3610 = _T_3589 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21863.4]
  assign _T_3611 = _T_3609 | _T_3610; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21864.4]
  assign _T_3613 = _T_3611 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21866.4]
  assign _T_3614 = _T_3613 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21867.4]
  assign _T_3625 = _T_2442 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21884.4]
  assign _T_3626 = _T_2702 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21885.4]
  assign _T_3628 = _T_3626 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21887.4]
  assign _T_3630 = _T_3620 + _T_3625; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21889.4]
  assign _T_3631 = _T_3630 - _T_3628; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21890.4]
  assign _T_3632 = $unsigned(_T_3631); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21891.4]
  assign _T_3633 = _T_3632[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21892.4]
  assign _T_3634 = _T_3628 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21894.4]
  assign _T_3636 = _T_3634 | _T_3620; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21896.4]
  assign _T_3638 = _T_3636 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21898.4]
  assign _T_3639 = _T_3638 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21899.4]
  assign _T_3640 = _T_3625 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21904.4]
  assign _T_3641 = _T_3620 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21905.4]
  assign _T_3642 = _T_3640 | _T_3641; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21906.4]
  assign _T_3644 = _T_3642 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21908.4]
  assign _T_3645 = _T_3644 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21909.4]
  assign _T_3656 = _T_2443 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21926.4]
  assign _T_3657 = _T_2703 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21927.4]
  assign _T_3659 = _T_3657 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21929.4]
  assign _T_3661 = _T_3651 + _T_3656; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21931.4]
  assign _T_3662 = _T_3661 - _T_3659; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21932.4]
  assign _T_3663 = $unsigned(_T_3662); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21933.4]
  assign _T_3664 = _T_3663[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21934.4]
  assign _T_3665 = _T_3659 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21936.4]
  assign _T_3667 = _T_3665 | _T_3651; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21938.4]
  assign _T_3669 = _T_3667 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21940.4]
  assign _T_3670 = _T_3669 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21941.4]
  assign _T_3671 = _T_3656 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21946.4]
  assign _T_3672 = _T_3651 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21947.4]
  assign _T_3673 = _T_3671 | _T_3672; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21948.4]
  assign _T_3675 = _T_3673 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21950.4]
  assign _T_3676 = _T_3675 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21951.4]
  assign _T_3687 = _T_2444 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@21968.4]
  assign _T_3688 = _T_2704 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@21969.4]
  assign _T_3690 = _T_3688 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@21971.4]
  assign _T_3692 = _T_3682 + _T_3687; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@21973.4]
  assign _T_3693 = _T_3692 - _T_3690; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21974.4]
  assign _T_3694 = $unsigned(_T_3693); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21975.4]
  assign _T_3695 = _T_3694[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@21976.4]
  assign _T_3696 = _T_3690 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@21978.4]
  assign _T_3698 = _T_3696 | _T_3682; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@21980.4]
  assign _T_3700 = _T_3698 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21982.4]
  assign _T_3701 = _T_3700 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21983.4]
  assign _T_3702 = _T_3687 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@21988.4]
  assign _T_3703 = _T_3682 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@21989.4]
  assign _T_3704 = _T_3702 | _T_3703; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@21990.4]
  assign _T_3706 = _T_3704 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21992.4]
  assign _T_3707 = _T_3706 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21993.4]
  assign _T_3718 = _T_2445 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22010.4]
  assign _T_3719 = _T_2705 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22011.4]
  assign _T_3721 = _T_3719 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22013.4]
  assign _T_3723 = _T_3713 + _T_3718; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22015.4]
  assign _T_3724 = _T_3723 - _T_3721; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22016.4]
  assign _T_3725 = $unsigned(_T_3724); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22017.4]
  assign _T_3726 = _T_3725[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22018.4]
  assign _T_3727 = _T_3721 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22020.4]
  assign _T_3729 = _T_3727 | _T_3713; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22022.4]
  assign _T_3731 = _T_3729 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22024.4]
  assign _T_3732 = _T_3731 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22025.4]
  assign _T_3733 = _T_3718 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22030.4]
  assign _T_3734 = _T_3713 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22031.4]
  assign _T_3735 = _T_3733 | _T_3734; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22032.4]
  assign _T_3737 = _T_3735 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22034.4]
  assign _T_3738 = _T_3737 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22035.4]
  assign _T_3749 = _T_2446 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22052.4]
  assign _T_3750 = _T_2706 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22053.4]
  assign _T_3752 = _T_3750 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22055.4]
  assign _T_3754 = _T_3744 + _T_3749; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22057.4]
  assign _T_3755 = _T_3754 - _T_3752; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22058.4]
  assign _T_3756 = $unsigned(_T_3755); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22059.4]
  assign _T_3757 = _T_3756[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22060.4]
  assign _T_3758 = _T_3752 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22062.4]
  assign _T_3760 = _T_3758 | _T_3744; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22064.4]
  assign _T_3762 = _T_3760 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22066.4]
  assign _T_3763 = _T_3762 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22067.4]
  assign _T_3764 = _T_3749 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22072.4]
  assign _T_3765 = _T_3744 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22073.4]
  assign _T_3766 = _T_3764 | _T_3765; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22074.4]
  assign _T_3768 = _T_3766 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22076.4]
  assign _T_3769 = _T_3768 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22077.4]
  assign _T_3780 = _T_2447 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22094.4]
  assign _T_3781 = _T_2707 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22095.4]
  assign _T_3783 = _T_3781 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22097.4]
  assign _T_3785 = _T_3775 + _T_3780; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22099.4]
  assign _T_3786 = _T_3785 - _T_3783; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22100.4]
  assign _T_3787 = $unsigned(_T_3786); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22101.4]
  assign _T_3788 = _T_3787[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22102.4]
  assign _T_3789 = _T_3783 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22104.4]
  assign _T_3791 = _T_3789 | _T_3775; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22106.4]
  assign _T_3793 = _T_3791 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22108.4]
  assign _T_3794 = _T_3793 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22109.4]
  assign _T_3795 = _T_3780 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22114.4]
  assign _T_3796 = _T_3775 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22115.4]
  assign _T_3797 = _T_3795 | _T_3796; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22116.4]
  assign _T_3799 = _T_3797 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22118.4]
  assign _T_3800 = _T_3799 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22119.4]
  assign _T_3811 = _T_2448 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22136.4]
  assign _T_3812 = _T_2708 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22137.4]
  assign _T_3814 = _T_3812 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22139.4]
  assign _T_3816 = _T_3806 + _T_3811; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22141.4]
  assign _T_3817 = _T_3816 - _T_3814; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22142.4]
  assign _T_3818 = $unsigned(_T_3817); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22143.4]
  assign _T_3819 = _T_3818[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22144.4]
  assign _T_3820 = _T_3814 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22146.4]
  assign _T_3822 = _T_3820 | _T_3806; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22148.4]
  assign _T_3824 = _T_3822 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22150.4]
  assign _T_3825 = _T_3824 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22151.4]
  assign _T_3826 = _T_3811 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22156.4]
  assign _T_3827 = _T_3806 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22157.4]
  assign _T_3828 = _T_3826 | _T_3827; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22158.4]
  assign _T_3830 = _T_3828 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22160.4]
  assign _T_3831 = _T_3830 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22161.4]
  assign _T_3842 = _T_2449 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22178.4]
  assign _T_3843 = _T_2709 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22179.4]
  assign _T_3845 = _T_3843 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22181.4]
  assign _T_3847 = _T_3837 + _T_3842; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22183.4]
  assign _T_3848 = _T_3847 - _T_3845; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22184.4]
  assign _T_3849 = $unsigned(_T_3848); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22185.4]
  assign _T_3850 = _T_3849[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22186.4]
  assign _T_3851 = _T_3845 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22188.4]
  assign _T_3853 = _T_3851 | _T_3837; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22190.4]
  assign _T_3855 = _T_3853 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22192.4]
  assign _T_3856 = _T_3855 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22193.4]
  assign _T_3857 = _T_3842 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22198.4]
  assign _T_3858 = _T_3837 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22199.4]
  assign _T_3859 = _T_3857 | _T_3858; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22200.4]
  assign _T_3861 = _T_3859 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22202.4]
  assign _T_3862 = _T_3861 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22203.4]
  assign _T_3873 = _T_2450 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22220.4]
  assign _T_3874 = _T_2710 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22221.4]
  assign _T_3876 = _T_3874 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22223.4]
  assign _T_3878 = _T_3868 + _T_3873; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22225.4]
  assign _T_3879 = _T_3878 - _T_3876; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22226.4]
  assign _T_3880 = $unsigned(_T_3879); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22227.4]
  assign _T_3881 = _T_3880[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22228.4]
  assign _T_3882 = _T_3876 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22230.4]
  assign _T_3884 = _T_3882 | _T_3868; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22232.4]
  assign _T_3886 = _T_3884 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22234.4]
  assign _T_3887 = _T_3886 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22235.4]
  assign _T_3888 = _T_3873 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22240.4]
  assign _T_3889 = _T_3868 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22241.4]
  assign _T_3890 = _T_3888 | _T_3889; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22242.4]
  assign _T_3892 = _T_3890 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22244.4]
  assign _T_3893 = _T_3892 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22245.4]
  assign _T_3904 = _T_2451 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22262.4]
  assign _T_3905 = _T_2711 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22263.4]
  assign _T_3907 = _T_3905 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22265.4]
  assign _T_3909 = _T_3899 + _T_3904; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22267.4]
  assign _T_3910 = _T_3909 - _T_3907; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22268.4]
  assign _T_3911 = $unsigned(_T_3910); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22269.4]
  assign _T_3912 = _T_3911[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22270.4]
  assign _T_3913 = _T_3907 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22272.4]
  assign _T_3915 = _T_3913 | _T_3899; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22274.4]
  assign _T_3917 = _T_3915 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22276.4]
  assign _T_3918 = _T_3917 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22277.4]
  assign _T_3919 = _T_3904 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22282.4]
  assign _T_3920 = _T_3899 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22283.4]
  assign _T_3921 = _T_3919 | _T_3920; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22284.4]
  assign _T_3923 = _T_3921 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22286.4]
  assign _T_3924 = _T_3923 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22287.4]
  assign _T_3935 = _T_2452 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22304.4]
  assign _T_3936 = _T_2712 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22305.4]
  assign _T_3938 = _T_3936 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22307.4]
  assign _T_3940 = _T_3930 + _T_3935; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22309.4]
  assign _T_3941 = _T_3940 - _T_3938; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22310.4]
  assign _T_3942 = $unsigned(_T_3941); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22311.4]
  assign _T_3943 = _T_3942[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22312.4]
  assign _T_3944 = _T_3938 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22314.4]
  assign _T_3946 = _T_3944 | _T_3930; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22316.4]
  assign _T_3948 = _T_3946 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22318.4]
  assign _T_3949 = _T_3948 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22319.4]
  assign _T_3950 = _T_3935 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22324.4]
  assign _T_3951 = _T_3930 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22325.4]
  assign _T_3952 = _T_3950 | _T_3951; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22326.4]
  assign _T_3954 = _T_3952 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22328.4]
  assign _T_3955 = _T_3954 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22329.4]
  assign _T_3966 = _T_2453 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22346.4]
  assign _T_3967 = _T_2713 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22347.4]
  assign _T_3969 = _T_3967 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22349.4]
  assign _T_3971 = _T_3961 + _T_3966; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22351.4]
  assign _T_3972 = _T_3971 - _T_3969; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22352.4]
  assign _T_3973 = $unsigned(_T_3972); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22353.4]
  assign _T_3974 = _T_3973[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22354.4]
  assign _T_3975 = _T_3969 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22356.4]
  assign _T_3977 = _T_3975 | _T_3961; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22358.4]
  assign _T_3979 = _T_3977 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22360.4]
  assign _T_3980 = _T_3979 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22361.4]
  assign _T_3981 = _T_3966 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22366.4]
  assign _T_3982 = _T_3961 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22367.4]
  assign _T_3983 = _T_3981 | _T_3982; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22368.4]
  assign _T_3985 = _T_3983 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22370.4]
  assign _T_3986 = _T_3985 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22371.4]
  assign _T_3997 = _T_2454 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22388.4]
  assign _T_3998 = _T_2714 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22389.4]
  assign _T_4000 = _T_3998 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22391.4]
  assign _T_4002 = _T_3992 + _T_3997; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22393.4]
  assign _T_4003 = _T_4002 - _T_4000; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22394.4]
  assign _T_4004 = $unsigned(_T_4003); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22395.4]
  assign _T_4005 = _T_4004[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22396.4]
  assign _T_4006 = _T_4000 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22398.4]
  assign _T_4008 = _T_4006 | _T_3992; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22400.4]
  assign _T_4010 = _T_4008 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22402.4]
  assign _T_4011 = _T_4010 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22403.4]
  assign _T_4012 = _T_3997 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22408.4]
  assign _T_4013 = _T_3992 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22409.4]
  assign _T_4014 = _T_4012 | _T_4013; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22410.4]
  assign _T_4016 = _T_4014 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22412.4]
  assign _T_4017 = _T_4016 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22413.4]
  assign _T_4028 = _T_2455 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22430.4]
  assign _T_4029 = _T_2715 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22431.4]
  assign _T_4031 = _T_4029 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22433.4]
  assign _T_4033 = _T_4023 + _T_4028; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22435.4]
  assign _T_4034 = _T_4033 - _T_4031; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22436.4]
  assign _T_4035 = $unsigned(_T_4034); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22437.4]
  assign _T_4036 = _T_4035[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22438.4]
  assign _T_4037 = _T_4031 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22440.4]
  assign _T_4039 = _T_4037 | _T_4023; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22442.4]
  assign _T_4041 = _T_4039 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22444.4]
  assign _T_4042 = _T_4041 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22445.4]
  assign _T_4043 = _T_4028 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22450.4]
  assign _T_4044 = _T_4023 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22451.4]
  assign _T_4045 = _T_4043 | _T_4044; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22452.4]
  assign _T_4047 = _T_4045 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22454.4]
  assign _T_4048 = _T_4047 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22455.4]
  assign _T_4059 = _T_2456 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22472.4]
  assign _T_4060 = _T_2716 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22473.4]
  assign _T_4062 = _T_4060 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22475.4]
  assign _T_4064 = _T_4054 + _T_4059; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22477.4]
  assign _T_4065 = _T_4064 - _T_4062; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22478.4]
  assign _T_4066 = $unsigned(_T_4065); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22479.4]
  assign _T_4067 = _T_4066[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22480.4]
  assign _T_4068 = _T_4062 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22482.4]
  assign _T_4070 = _T_4068 | _T_4054; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22484.4]
  assign _T_4072 = _T_4070 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22486.4]
  assign _T_4073 = _T_4072 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22487.4]
  assign _T_4074 = _T_4059 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22492.4]
  assign _T_4075 = _T_4054 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22493.4]
  assign _T_4076 = _T_4074 | _T_4075; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22494.4]
  assign _T_4078 = _T_4076 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22496.4]
  assign _T_4079 = _T_4078 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22497.4]
  assign _T_4090 = _T_2457 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22514.4]
  assign _T_4091 = _T_2717 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22515.4]
  assign _T_4093 = _T_4091 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22517.4]
  assign _T_4095 = _T_4085 + _T_4090; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22519.4]
  assign _T_4096 = _T_4095 - _T_4093; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22520.4]
  assign _T_4097 = $unsigned(_T_4096); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22521.4]
  assign _T_4098 = _T_4097[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22522.4]
  assign _T_4099 = _T_4093 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22524.4]
  assign _T_4101 = _T_4099 | _T_4085; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22526.4]
  assign _T_4103 = _T_4101 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22528.4]
  assign _T_4104 = _T_4103 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22529.4]
  assign _T_4105 = _T_4090 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22534.4]
  assign _T_4106 = _T_4085 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22535.4]
  assign _T_4107 = _T_4105 | _T_4106; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22536.4]
  assign _T_4109 = _T_4107 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22538.4]
  assign _T_4110 = _T_4109 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22539.4]
  assign _T_4121 = _T_2458 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22556.4]
  assign _T_4122 = _T_2718 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22557.4]
  assign _T_4124 = _T_4122 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22559.4]
  assign _T_4126 = _T_4116 + _T_4121; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22561.4]
  assign _T_4127 = _T_4126 - _T_4124; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22562.4]
  assign _T_4128 = $unsigned(_T_4127); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22563.4]
  assign _T_4129 = _T_4128[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22564.4]
  assign _T_4130 = _T_4124 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22566.4]
  assign _T_4132 = _T_4130 | _T_4116; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22568.4]
  assign _T_4134 = _T_4132 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22570.4]
  assign _T_4135 = _T_4134 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22571.4]
  assign _T_4136 = _T_4121 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22576.4]
  assign _T_4137 = _T_4116 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22577.4]
  assign _T_4138 = _T_4136 | _T_4137; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22578.4]
  assign _T_4140 = _T_4138 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22580.4]
  assign _T_4141 = _T_4140 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22581.4]
  assign _T_4152 = _T_2459 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22598.4]
  assign _T_4153 = _T_2719 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22599.4]
  assign _T_4155 = _T_4153 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22601.4]
  assign _T_4157 = _T_4147 + _T_4152; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22603.4]
  assign _T_4158 = _T_4157 - _T_4155; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22604.4]
  assign _T_4159 = $unsigned(_T_4158); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22605.4]
  assign _T_4160 = _T_4159[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22606.4]
  assign _T_4161 = _T_4155 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22608.4]
  assign _T_4163 = _T_4161 | _T_4147; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22610.4]
  assign _T_4165 = _T_4163 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22612.4]
  assign _T_4166 = _T_4165 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22613.4]
  assign _T_4167 = _T_4152 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22618.4]
  assign _T_4168 = _T_4147 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22619.4]
  assign _T_4169 = _T_4167 | _T_4168; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22620.4]
  assign _T_4171 = _T_4169 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22622.4]
  assign _T_4172 = _T_4171 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22623.4]
  assign _T_4183 = _T_2460 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22640.4]
  assign _T_4184 = _T_2720 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22641.4]
  assign _T_4186 = _T_4184 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22643.4]
  assign _T_4188 = _T_4178 + _T_4183; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22645.4]
  assign _T_4189 = _T_4188 - _T_4186; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22646.4]
  assign _T_4190 = $unsigned(_T_4189); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22647.4]
  assign _T_4191 = _T_4190[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22648.4]
  assign _T_4192 = _T_4186 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22650.4]
  assign _T_4194 = _T_4192 | _T_4178; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22652.4]
  assign _T_4196 = _T_4194 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22654.4]
  assign _T_4197 = _T_4196 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22655.4]
  assign _T_4198 = _T_4183 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22660.4]
  assign _T_4199 = _T_4178 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22661.4]
  assign _T_4200 = _T_4198 | _T_4199; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22662.4]
  assign _T_4202 = _T_4200 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22664.4]
  assign _T_4203 = _T_4202 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22665.4]
  assign _T_4214 = _T_2461 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22682.4]
  assign _T_4215 = _T_2721 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22683.4]
  assign _T_4217 = _T_4215 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22685.4]
  assign _T_4219 = _T_4209 + _T_4214; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22687.4]
  assign _T_4220 = _T_4219 - _T_4217; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22688.4]
  assign _T_4221 = $unsigned(_T_4220); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22689.4]
  assign _T_4222 = _T_4221[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22690.4]
  assign _T_4223 = _T_4217 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22692.4]
  assign _T_4225 = _T_4223 | _T_4209; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22694.4]
  assign _T_4227 = _T_4225 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22696.4]
  assign _T_4228 = _T_4227 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22697.4]
  assign _T_4229 = _T_4214 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22702.4]
  assign _T_4230 = _T_4209 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22703.4]
  assign _T_4231 = _T_4229 | _T_4230; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22704.4]
  assign _T_4233 = _T_4231 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22706.4]
  assign _T_4234 = _T_4233 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22707.4]
  assign _T_4245 = _T_2462 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22724.4]
  assign _T_4246 = _T_2722 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22725.4]
  assign _T_4248 = _T_4246 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22727.4]
  assign _T_4250 = _T_4240 + _T_4245; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22729.4]
  assign _T_4251 = _T_4250 - _T_4248; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22730.4]
  assign _T_4252 = $unsigned(_T_4251); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22731.4]
  assign _T_4253 = _T_4252[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22732.4]
  assign _T_4254 = _T_4248 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22734.4]
  assign _T_4256 = _T_4254 | _T_4240; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22736.4]
  assign _T_4258 = _T_4256 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22738.4]
  assign _T_4259 = _T_4258 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22739.4]
  assign _T_4260 = _T_4245 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22744.4]
  assign _T_4261 = _T_4240 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22745.4]
  assign _T_4262 = _T_4260 | _T_4261; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22746.4]
  assign _T_4264 = _T_4262 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22748.4]
  assign _T_4265 = _T_4264 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22749.4]
  assign _T_4276 = _T_2463 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22766.4]
  assign _T_4277 = _T_2723 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22767.4]
  assign _T_4279 = _T_4277 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22769.4]
  assign _T_4281 = _T_4271 + _T_4276; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22771.4]
  assign _T_4282 = _T_4281 - _T_4279; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22772.4]
  assign _T_4283 = $unsigned(_T_4282); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22773.4]
  assign _T_4284 = _T_4283[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22774.4]
  assign _T_4285 = _T_4279 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22776.4]
  assign _T_4287 = _T_4285 | _T_4271; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22778.4]
  assign _T_4289 = _T_4287 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22780.4]
  assign _T_4290 = _T_4289 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22781.4]
  assign _T_4291 = _T_4276 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22786.4]
  assign _T_4292 = _T_4271 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22787.4]
  assign _T_4293 = _T_4291 | _T_4292; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22788.4]
  assign _T_4295 = _T_4293 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22790.4]
  assign _T_4296 = _T_4295 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22791.4]
  assign _T_4307 = _T_2464 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22808.4]
  assign _T_4308 = _T_2724 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22809.4]
  assign _T_4310 = _T_4308 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22811.4]
  assign _T_4312 = _T_4302 + _T_4307; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22813.4]
  assign _T_4313 = _T_4312 - _T_4310; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22814.4]
  assign _T_4314 = $unsigned(_T_4313); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22815.4]
  assign _T_4315 = _T_4314[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22816.4]
  assign _T_4316 = _T_4310 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22818.4]
  assign _T_4318 = _T_4316 | _T_4302; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22820.4]
  assign _T_4320 = _T_4318 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22822.4]
  assign _T_4321 = _T_4320 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22823.4]
  assign _T_4322 = _T_4307 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22828.4]
  assign _T_4323 = _T_4302 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22829.4]
  assign _T_4324 = _T_4322 | _T_4323; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22830.4]
  assign _T_4326 = _T_4324 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22832.4]
  assign _T_4327 = _T_4326 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22833.4]
  assign _T_4338 = _T_2465 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22850.4]
  assign _T_4339 = _T_2725 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22851.4]
  assign _T_4341 = _T_4339 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22853.4]
  assign _T_4343 = _T_4333 + _T_4338; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22855.4]
  assign _T_4344 = _T_4343 - _T_4341; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22856.4]
  assign _T_4345 = $unsigned(_T_4344); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22857.4]
  assign _T_4346 = _T_4345[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22858.4]
  assign _T_4347 = _T_4341 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22860.4]
  assign _T_4349 = _T_4347 | _T_4333; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22862.4]
  assign _T_4351 = _T_4349 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22864.4]
  assign _T_4352 = _T_4351 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22865.4]
  assign _T_4353 = _T_4338 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22870.4]
  assign _T_4354 = _T_4333 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22871.4]
  assign _T_4355 = _T_4353 | _T_4354; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22872.4]
  assign _T_4357 = _T_4355 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22874.4]
  assign _T_4358 = _T_4357 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22875.4]
  assign _T_4369 = _T_2466 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22892.4]
  assign _T_4370 = _T_2726 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22893.4]
  assign _T_4372 = _T_4370 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22895.4]
  assign _T_4374 = _T_4364 + _T_4369; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22897.4]
  assign _T_4375 = _T_4374 - _T_4372; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22898.4]
  assign _T_4376 = $unsigned(_T_4375); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22899.4]
  assign _T_4377 = _T_4376[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22900.4]
  assign _T_4378 = _T_4372 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22902.4]
  assign _T_4380 = _T_4378 | _T_4364; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22904.4]
  assign _T_4382 = _T_4380 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22906.4]
  assign _T_4383 = _T_4382 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22907.4]
  assign _T_4384 = _T_4369 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22912.4]
  assign _T_4385 = _T_4364 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22913.4]
  assign _T_4386 = _T_4384 | _T_4385; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22914.4]
  assign _T_4388 = _T_4386 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22916.4]
  assign _T_4389 = _T_4388 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22917.4]
  assign _T_4400 = _T_2467 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22934.4]
  assign _T_4401 = _T_2727 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22935.4]
  assign _T_4403 = _T_4401 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22937.4]
  assign _T_4405 = _T_4395 + _T_4400; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22939.4]
  assign _T_4406 = _T_4405 - _T_4403; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22940.4]
  assign _T_4407 = $unsigned(_T_4406); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22941.4]
  assign _T_4408 = _T_4407[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22942.4]
  assign _T_4409 = _T_4403 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22944.4]
  assign _T_4411 = _T_4409 | _T_4395; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22946.4]
  assign _T_4413 = _T_4411 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22948.4]
  assign _T_4414 = _T_4413 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22949.4]
  assign _T_4415 = _T_4400 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22954.4]
  assign _T_4416 = _T_4395 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22955.4]
  assign _T_4417 = _T_4415 | _T_4416; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22956.4]
  assign _T_4419 = _T_4417 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22958.4]
  assign _T_4420 = _T_4419 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22959.4]
  assign _T_4431 = _T_2468 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@22976.4]
  assign _T_4432 = _T_2728 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@22977.4]
  assign _T_4434 = _T_4432 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@22979.4]
  assign _T_4436 = _T_4426 + _T_4431; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@22981.4]
  assign _T_4437 = _T_4436 - _T_4434; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22982.4]
  assign _T_4438 = $unsigned(_T_4437); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22983.4]
  assign _T_4439 = _T_4438[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@22984.4]
  assign _T_4440 = _T_4434 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@22986.4]
  assign _T_4442 = _T_4440 | _T_4426; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@22988.4]
  assign _T_4444 = _T_4442 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22990.4]
  assign _T_4445 = _T_4444 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22991.4]
  assign _T_4446 = _T_4431 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@22996.4]
  assign _T_4447 = _T_4426 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@22997.4]
  assign _T_4448 = _T_4446 | _T_4447; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@22998.4]
  assign _T_4450 = _T_4448 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23000.4]
  assign _T_4451 = _T_4450 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23001.4]
  assign _T_4462 = _T_2469 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23018.4]
  assign _T_4463 = _T_2729 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23019.4]
  assign _T_4465 = _T_4463 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23021.4]
  assign _T_4467 = _T_4457 + _T_4462; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23023.4]
  assign _T_4468 = _T_4467 - _T_4465; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23024.4]
  assign _T_4469 = $unsigned(_T_4468); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23025.4]
  assign _T_4470 = _T_4469[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23026.4]
  assign _T_4471 = _T_4465 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23028.4]
  assign _T_4473 = _T_4471 | _T_4457; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23030.4]
  assign _T_4475 = _T_4473 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23032.4]
  assign _T_4476 = _T_4475 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23033.4]
  assign _T_4477 = _T_4462 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23038.4]
  assign _T_4478 = _T_4457 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23039.4]
  assign _T_4479 = _T_4477 | _T_4478; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23040.4]
  assign _T_4481 = _T_4479 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23042.4]
  assign _T_4482 = _T_4481 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23043.4]
  assign _T_4493 = _T_2470 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23060.4]
  assign _T_4494 = _T_2730 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23061.4]
  assign _T_4496 = _T_4494 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23063.4]
  assign _T_4498 = _T_4488 + _T_4493; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23065.4]
  assign _T_4499 = _T_4498 - _T_4496; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23066.4]
  assign _T_4500 = $unsigned(_T_4499); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23067.4]
  assign _T_4501 = _T_4500[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23068.4]
  assign _T_4502 = _T_4496 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23070.4]
  assign _T_4504 = _T_4502 | _T_4488; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23072.4]
  assign _T_4506 = _T_4504 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23074.4]
  assign _T_4507 = _T_4506 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23075.4]
  assign _T_4508 = _T_4493 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23080.4]
  assign _T_4509 = _T_4488 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23081.4]
  assign _T_4510 = _T_4508 | _T_4509; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23082.4]
  assign _T_4512 = _T_4510 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23084.4]
  assign _T_4513 = _T_4512 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23085.4]
  assign _T_4524 = _T_2471 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23102.4]
  assign _T_4525 = _T_2731 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23103.4]
  assign _T_4527 = _T_4525 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23105.4]
  assign _T_4529 = _T_4519 + _T_4524; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23107.4]
  assign _T_4530 = _T_4529 - _T_4527; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23108.4]
  assign _T_4531 = $unsigned(_T_4530); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23109.4]
  assign _T_4532 = _T_4531[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23110.4]
  assign _T_4533 = _T_4527 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23112.4]
  assign _T_4535 = _T_4533 | _T_4519; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23114.4]
  assign _T_4537 = _T_4535 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23116.4]
  assign _T_4538 = _T_4537 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23117.4]
  assign _T_4539 = _T_4524 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23122.4]
  assign _T_4540 = _T_4519 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23123.4]
  assign _T_4541 = _T_4539 | _T_4540; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23124.4]
  assign _T_4543 = _T_4541 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23126.4]
  assign _T_4544 = _T_4543 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23127.4]
  assign _T_4555 = _T_2472 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23144.4]
  assign _T_4556 = _T_2732 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23145.4]
  assign _T_4558 = _T_4556 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23147.4]
  assign _T_4560 = _T_4550 + _T_4555; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23149.4]
  assign _T_4561 = _T_4560 - _T_4558; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23150.4]
  assign _T_4562 = $unsigned(_T_4561); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23151.4]
  assign _T_4563 = _T_4562[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23152.4]
  assign _T_4564 = _T_4558 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23154.4]
  assign _T_4566 = _T_4564 | _T_4550; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23156.4]
  assign _T_4568 = _T_4566 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23158.4]
  assign _T_4569 = _T_4568 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23159.4]
  assign _T_4570 = _T_4555 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23164.4]
  assign _T_4571 = _T_4550 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23165.4]
  assign _T_4572 = _T_4570 | _T_4571; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23166.4]
  assign _T_4574 = _T_4572 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23168.4]
  assign _T_4575 = _T_4574 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23169.4]
  assign _T_4586 = _T_2473 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23186.4]
  assign _T_4587 = _T_2733 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23187.4]
  assign _T_4589 = _T_4587 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23189.4]
  assign _T_4591 = _T_4581 + _T_4586; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23191.4]
  assign _T_4592 = _T_4591 - _T_4589; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23192.4]
  assign _T_4593 = $unsigned(_T_4592); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23193.4]
  assign _T_4594 = _T_4593[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23194.4]
  assign _T_4595 = _T_4589 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23196.4]
  assign _T_4597 = _T_4595 | _T_4581; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23198.4]
  assign _T_4599 = _T_4597 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23200.4]
  assign _T_4600 = _T_4599 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23201.4]
  assign _T_4601 = _T_4586 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23206.4]
  assign _T_4602 = _T_4581 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23207.4]
  assign _T_4603 = _T_4601 | _T_4602; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23208.4]
  assign _T_4605 = _T_4603 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23210.4]
  assign _T_4606 = _T_4605 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23211.4]
  assign _T_4617 = _T_2474 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23228.4]
  assign _T_4618 = _T_2734 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23229.4]
  assign _T_4620 = _T_4618 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23231.4]
  assign _T_4622 = _T_4612 + _T_4617; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23233.4]
  assign _T_4623 = _T_4622 - _T_4620; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23234.4]
  assign _T_4624 = $unsigned(_T_4623); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23235.4]
  assign _T_4625 = _T_4624[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23236.4]
  assign _T_4626 = _T_4620 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23238.4]
  assign _T_4628 = _T_4626 | _T_4612; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23240.4]
  assign _T_4630 = _T_4628 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23242.4]
  assign _T_4631 = _T_4630 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23243.4]
  assign _T_4632 = _T_4617 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23248.4]
  assign _T_4633 = _T_4612 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23249.4]
  assign _T_4634 = _T_4632 | _T_4633; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23250.4]
  assign _T_4636 = _T_4634 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23252.4]
  assign _T_4637 = _T_4636 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23253.4]
  assign _T_4648 = _T_2475 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23270.4]
  assign _T_4649 = _T_2735 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23271.4]
  assign _T_4651 = _T_4649 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23273.4]
  assign _T_4653 = _T_4643 + _T_4648; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23275.4]
  assign _T_4654 = _T_4653 - _T_4651; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23276.4]
  assign _T_4655 = $unsigned(_T_4654); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23277.4]
  assign _T_4656 = _T_4655[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23278.4]
  assign _T_4657 = _T_4651 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23280.4]
  assign _T_4659 = _T_4657 | _T_4643; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23282.4]
  assign _T_4661 = _T_4659 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23284.4]
  assign _T_4662 = _T_4661 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23285.4]
  assign _T_4663 = _T_4648 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23290.4]
  assign _T_4664 = _T_4643 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23291.4]
  assign _T_4665 = _T_4663 | _T_4664; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23292.4]
  assign _T_4667 = _T_4665 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23294.4]
  assign _T_4668 = _T_4667 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23295.4]
  assign _T_4679 = _T_2476 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23312.4]
  assign _T_4680 = _T_2736 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23313.4]
  assign _T_4682 = _T_4680 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23315.4]
  assign _T_4684 = _T_4674 + _T_4679; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23317.4]
  assign _T_4685 = _T_4684 - _T_4682; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23318.4]
  assign _T_4686 = $unsigned(_T_4685); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23319.4]
  assign _T_4687 = _T_4686[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23320.4]
  assign _T_4688 = _T_4682 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23322.4]
  assign _T_4690 = _T_4688 | _T_4674; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23324.4]
  assign _T_4692 = _T_4690 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23326.4]
  assign _T_4693 = _T_4692 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23327.4]
  assign _T_4694 = _T_4679 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23332.4]
  assign _T_4695 = _T_4674 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23333.4]
  assign _T_4696 = _T_4694 | _T_4695; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23334.4]
  assign _T_4698 = _T_4696 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23336.4]
  assign _T_4699 = _T_4698 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23337.4]
  assign _T_4710 = _T_2477 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23354.4]
  assign _T_4711 = _T_2737 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23355.4]
  assign _T_4713 = _T_4711 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23357.4]
  assign _T_4715 = _T_4705 + _T_4710; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23359.4]
  assign _T_4716 = _T_4715 - _T_4713; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23360.4]
  assign _T_4717 = $unsigned(_T_4716); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23361.4]
  assign _T_4718 = _T_4717[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23362.4]
  assign _T_4719 = _T_4713 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23364.4]
  assign _T_4721 = _T_4719 | _T_4705; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23366.4]
  assign _T_4723 = _T_4721 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23368.4]
  assign _T_4724 = _T_4723 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23369.4]
  assign _T_4725 = _T_4710 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23374.4]
  assign _T_4726 = _T_4705 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23375.4]
  assign _T_4727 = _T_4725 | _T_4726; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23376.4]
  assign _T_4729 = _T_4727 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23378.4]
  assign _T_4730 = _T_4729 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23379.4]
  assign _T_4741 = _T_2478 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23396.4]
  assign _T_4742 = _T_2738 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23397.4]
  assign _T_4744 = _T_4742 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23399.4]
  assign _T_4746 = _T_4736 + _T_4741; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23401.4]
  assign _T_4747 = _T_4746 - _T_4744; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23402.4]
  assign _T_4748 = $unsigned(_T_4747); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23403.4]
  assign _T_4749 = _T_4748[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23404.4]
  assign _T_4750 = _T_4744 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23406.4]
  assign _T_4752 = _T_4750 | _T_4736; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23408.4]
  assign _T_4754 = _T_4752 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23410.4]
  assign _T_4755 = _T_4754 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23411.4]
  assign _T_4756 = _T_4741 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23416.4]
  assign _T_4757 = _T_4736 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23417.4]
  assign _T_4758 = _T_4756 | _T_4757; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23418.4]
  assign _T_4760 = _T_4758 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23420.4]
  assign _T_4761 = _T_4760 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23421.4]
  assign _T_4772 = _T_2479 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23438.4]
  assign _T_4773 = _T_2739 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23439.4]
  assign _T_4775 = _T_4773 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23441.4]
  assign _T_4777 = _T_4767 + _T_4772; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23443.4]
  assign _T_4778 = _T_4777 - _T_4775; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23444.4]
  assign _T_4779 = $unsigned(_T_4778); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23445.4]
  assign _T_4780 = _T_4779[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23446.4]
  assign _T_4781 = _T_4775 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23448.4]
  assign _T_4783 = _T_4781 | _T_4767; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23450.4]
  assign _T_4785 = _T_4783 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23452.4]
  assign _T_4786 = _T_4785 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23453.4]
  assign _T_4787 = _T_4772 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23458.4]
  assign _T_4788 = _T_4767 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23459.4]
  assign _T_4789 = _T_4787 | _T_4788; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23460.4]
  assign _T_4791 = _T_4789 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23462.4]
  assign _T_4792 = _T_4791 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23463.4]
  assign _T_4803 = _T_2480 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23480.4]
  assign _T_4804 = _T_2740 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23481.4]
  assign _T_4806 = _T_4804 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23483.4]
  assign _T_4808 = _T_4798 + _T_4803; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23485.4]
  assign _T_4809 = _T_4808 - _T_4806; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23486.4]
  assign _T_4810 = $unsigned(_T_4809); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23487.4]
  assign _T_4811 = _T_4810[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23488.4]
  assign _T_4812 = _T_4806 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23490.4]
  assign _T_4814 = _T_4812 | _T_4798; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23492.4]
  assign _T_4816 = _T_4814 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23494.4]
  assign _T_4817 = _T_4816 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23495.4]
  assign _T_4818 = _T_4803 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23500.4]
  assign _T_4819 = _T_4798 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23501.4]
  assign _T_4820 = _T_4818 | _T_4819; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23502.4]
  assign _T_4822 = _T_4820 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23504.4]
  assign _T_4823 = _T_4822 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23505.4]
  assign _T_4834 = _T_2481 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23522.4]
  assign _T_4835 = _T_2741 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23523.4]
  assign _T_4837 = _T_4835 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23525.4]
  assign _T_4839 = _T_4829 + _T_4834; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23527.4]
  assign _T_4840 = _T_4839 - _T_4837; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23528.4]
  assign _T_4841 = $unsigned(_T_4840); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23529.4]
  assign _T_4842 = _T_4841[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23530.4]
  assign _T_4843 = _T_4837 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23532.4]
  assign _T_4845 = _T_4843 | _T_4829; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23534.4]
  assign _T_4847 = _T_4845 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23536.4]
  assign _T_4848 = _T_4847 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23537.4]
  assign _T_4849 = _T_4834 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23542.4]
  assign _T_4850 = _T_4829 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23543.4]
  assign _T_4851 = _T_4849 | _T_4850; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23544.4]
  assign _T_4853 = _T_4851 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23546.4]
  assign _T_4854 = _T_4853 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23547.4]
  assign _T_4865 = _T_2482 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23564.4]
  assign _T_4866 = _T_2742 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23565.4]
  assign _T_4868 = _T_4866 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23567.4]
  assign _T_4870 = _T_4860 + _T_4865; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23569.4]
  assign _T_4871 = _T_4870 - _T_4868; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23570.4]
  assign _T_4872 = $unsigned(_T_4871); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23571.4]
  assign _T_4873 = _T_4872[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23572.4]
  assign _T_4874 = _T_4868 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23574.4]
  assign _T_4876 = _T_4874 | _T_4860; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23576.4]
  assign _T_4878 = _T_4876 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23578.4]
  assign _T_4879 = _T_4878 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23579.4]
  assign _T_4880 = _T_4865 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23584.4]
  assign _T_4881 = _T_4860 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23585.4]
  assign _T_4882 = _T_4880 | _T_4881; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23586.4]
  assign _T_4884 = _T_4882 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23588.4]
  assign _T_4885 = _T_4884 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23589.4]
  assign _T_4896 = _T_2483 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23606.4]
  assign _T_4897 = _T_2743 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23607.4]
  assign _T_4899 = _T_4897 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23609.4]
  assign _T_4901 = _T_4891 + _T_4896; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23611.4]
  assign _T_4902 = _T_4901 - _T_4899; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23612.4]
  assign _T_4903 = $unsigned(_T_4902); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23613.4]
  assign _T_4904 = _T_4903[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23614.4]
  assign _T_4905 = _T_4899 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23616.4]
  assign _T_4907 = _T_4905 | _T_4891; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23618.4]
  assign _T_4909 = _T_4907 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23620.4]
  assign _T_4910 = _T_4909 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23621.4]
  assign _T_4911 = _T_4896 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23626.4]
  assign _T_4912 = _T_4891 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23627.4]
  assign _T_4913 = _T_4911 | _T_4912; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23628.4]
  assign _T_4915 = _T_4913 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23630.4]
  assign _T_4916 = _T_4915 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23631.4]
  assign _T_4927 = _T_2484 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23648.4]
  assign _T_4928 = _T_2744 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23649.4]
  assign _T_4930 = _T_4928 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23651.4]
  assign _T_4932 = _T_4922 + _T_4927; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23653.4]
  assign _T_4933 = _T_4932 - _T_4930; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23654.4]
  assign _T_4934 = $unsigned(_T_4933); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23655.4]
  assign _T_4935 = _T_4934[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23656.4]
  assign _T_4936 = _T_4930 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23658.4]
  assign _T_4938 = _T_4936 | _T_4922; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23660.4]
  assign _T_4940 = _T_4938 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23662.4]
  assign _T_4941 = _T_4940 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23663.4]
  assign _T_4942 = _T_4927 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23668.4]
  assign _T_4943 = _T_4922 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23669.4]
  assign _T_4944 = _T_4942 | _T_4943; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23670.4]
  assign _T_4946 = _T_4944 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23672.4]
  assign _T_4947 = _T_4946 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23673.4]
  assign _T_4958 = _T_2485 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23690.4]
  assign _T_4959 = _T_2745 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23691.4]
  assign _T_4961 = _T_4959 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23693.4]
  assign _T_4963 = _T_4953 + _T_4958; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23695.4]
  assign _T_4964 = _T_4963 - _T_4961; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23696.4]
  assign _T_4965 = $unsigned(_T_4964); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23697.4]
  assign _T_4966 = _T_4965[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23698.4]
  assign _T_4967 = _T_4961 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23700.4]
  assign _T_4969 = _T_4967 | _T_4953; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23702.4]
  assign _T_4971 = _T_4969 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23704.4]
  assign _T_4972 = _T_4971 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23705.4]
  assign _T_4973 = _T_4958 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23710.4]
  assign _T_4974 = _T_4953 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23711.4]
  assign _T_4975 = _T_4973 | _T_4974; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23712.4]
  assign _T_4977 = _T_4975 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23714.4]
  assign _T_4978 = _T_4977 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23715.4]
  assign _T_4989 = _T_2486 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23732.4]
  assign _T_4990 = _T_2746 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23733.4]
  assign _T_4992 = _T_4990 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23735.4]
  assign _T_4994 = _T_4984 + _T_4989; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23737.4]
  assign _T_4995 = _T_4994 - _T_4992; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23738.4]
  assign _T_4996 = $unsigned(_T_4995); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23739.4]
  assign _T_4997 = _T_4996[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23740.4]
  assign _T_4998 = _T_4992 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23742.4]
  assign _T_5000 = _T_4998 | _T_4984; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23744.4]
  assign _T_5002 = _T_5000 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23746.4]
  assign _T_5003 = _T_5002 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23747.4]
  assign _T_5004 = _T_4989 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23752.4]
  assign _T_5005 = _T_4984 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23753.4]
  assign _T_5006 = _T_5004 | _T_5005; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23754.4]
  assign _T_5008 = _T_5006 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23756.4]
  assign _T_5009 = _T_5008 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23757.4]
  assign _T_5020 = _T_2487 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23774.4]
  assign _T_5021 = _T_2747 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23775.4]
  assign _T_5023 = _T_5021 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23777.4]
  assign _T_5025 = _T_5015 + _T_5020; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23779.4]
  assign _T_5026 = _T_5025 - _T_5023; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23780.4]
  assign _T_5027 = $unsigned(_T_5026); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23781.4]
  assign _T_5028 = _T_5027[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23782.4]
  assign _T_5029 = _T_5023 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23784.4]
  assign _T_5031 = _T_5029 | _T_5015; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23786.4]
  assign _T_5033 = _T_5031 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23788.4]
  assign _T_5034 = _T_5033 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23789.4]
  assign _T_5035 = _T_5020 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23794.4]
  assign _T_5036 = _T_5015 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23795.4]
  assign _T_5037 = _T_5035 | _T_5036; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23796.4]
  assign _T_5039 = _T_5037 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23798.4]
  assign _T_5040 = _T_5039 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23799.4]
  assign _T_5051 = _T_2488 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23816.4]
  assign _T_5052 = _T_2748 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23817.4]
  assign _T_5054 = _T_5052 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23819.4]
  assign _T_5056 = _T_5046 + _T_5051; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23821.4]
  assign _T_5057 = _T_5056 - _T_5054; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23822.4]
  assign _T_5058 = $unsigned(_T_5057); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23823.4]
  assign _T_5059 = _T_5058[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23824.4]
  assign _T_5060 = _T_5054 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23826.4]
  assign _T_5062 = _T_5060 | _T_5046; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23828.4]
  assign _T_5064 = _T_5062 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23830.4]
  assign _T_5065 = _T_5064 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23831.4]
  assign _T_5066 = _T_5051 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23836.4]
  assign _T_5067 = _T_5046 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23837.4]
  assign _T_5068 = _T_5066 | _T_5067; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23838.4]
  assign _T_5070 = _T_5068 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23840.4]
  assign _T_5071 = _T_5070 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23841.4]
  assign _T_5082 = _T_2489 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23858.4]
  assign _T_5083 = _T_2749 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23859.4]
  assign _T_5085 = _T_5083 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23861.4]
  assign _T_5087 = _T_5077 + _T_5082; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23863.4]
  assign _T_5088 = _T_5087 - _T_5085; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23864.4]
  assign _T_5089 = $unsigned(_T_5088); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23865.4]
  assign _T_5090 = _T_5089[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23866.4]
  assign _T_5091 = _T_5085 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23868.4]
  assign _T_5093 = _T_5091 | _T_5077; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23870.4]
  assign _T_5095 = _T_5093 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23872.4]
  assign _T_5096 = _T_5095 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23873.4]
  assign _T_5097 = _T_5082 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23878.4]
  assign _T_5098 = _T_5077 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23879.4]
  assign _T_5099 = _T_5097 | _T_5098; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23880.4]
  assign _T_5101 = _T_5099 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23882.4]
  assign _T_5102 = _T_5101 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23883.4]
  assign _T_5113 = _T_2490 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23900.4]
  assign _T_5114 = _T_2750 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23901.4]
  assign _T_5116 = _T_5114 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23903.4]
  assign _T_5118 = _T_5108 + _T_5113; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23905.4]
  assign _T_5119 = _T_5118 - _T_5116; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23906.4]
  assign _T_5120 = $unsigned(_T_5119); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23907.4]
  assign _T_5121 = _T_5120[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23908.4]
  assign _T_5122 = _T_5116 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23910.4]
  assign _T_5124 = _T_5122 | _T_5108; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23912.4]
  assign _T_5126 = _T_5124 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23914.4]
  assign _T_5127 = _T_5126 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23915.4]
  assign _T_5128 = _T_5113 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23920.4]
  assign _T_5129 = _T_5108 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23921.4]
  assign _T_5130 = _T_5128 | _T_5129; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23922.4]
  assign _T_5132 = _T_5130 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23924.4]
  assign _T_5133 = _T_5132 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23925.4]
  assign _T_5144 = _T_2491 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23942.4]
  assign _T_5145 = _T_2751 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23943.4]
  assign _T_5147 = _T_5145 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23945.4]
  assign _T_5149 = _T_5139 + _T_5144; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23947.4]
  assign _T_5150 = _T_5149 - _T_5147; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23948.4]
  assign _T_5151 = $unsigned(_T_5150); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23949.4]
  assign _T_5152 = _T_5151[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23950.4]
  assign _T_5153 = _T_5147 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23952.4]
  assign _T_5155 = _T_5153 | _T_5139; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23954.4]
  assign _T_5157 = _T_5155 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23956.4]
  assign _T_5158 = _T_5157 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23957.4]
  assign _T_5159 = _T_5144 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@23962.4]
  assign _T_5160 = _T_5139 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@23963.4]
  assign _T_5161 = _T_5159 | _T_5160; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@23964.4]
  assign _T_5163 = _T_5161 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23966.4]
  assign _T_5164 = _T_5163 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23967.4]
  assign _T_5175 = _T_2492 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@23984.4]
  assign _T_5176 = _T_2752 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@23985.4]
  assign _T_5178 = _T_5176 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@23987.4]
  assign _T_5180 = _T_5170 + _T_5175; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@23989.4]
  assign _T_5181 = _T_5180 - _T_5178; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23990.4]
  assign _T_5182 = $unsigned(_T_5181); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23991.4]
  assign _T_5183 = _T_5182[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@23992.4]
  assign _T_5184 = _T_5178 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@23994.4]
  assign _T_5186 = _T_5184 | _T_5170; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@23996.4]
  assign _T_5188 = _T_5186 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23998.4]
  assign _T_5189 = _T_5188 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23999.4]
  assign _T_5190 = _T_5175 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24004.4]
  assign _T_5191 = _T_5170 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24005.4]
  assign _T_5192 = _T_5190 | _T_5191; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24006.4]
  assign _T_5194 = _T_5192 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24008.4]
  assign _T_5195 = _T_5194 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24009.4]
  assign _T_5206 = _T_2493 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24026.4]
  assign _T_5207 = _T_2753 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24027.4]
  assign _T_5209 = _T_5207 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24029.4]
  assign _T_5211 = _T_5201 + _T_5206; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24031.4]
  assign _T_5212 = _T_5211 - _T_5209; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24032.4]
  assign _T_5213 = $unsigned(_T_5212); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24033.4]
  assign _T_5214 = _T_5213[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24034.4]
  assign _T_5215 = _T_5209 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24036.4]
  assign _T_5217 = _T_5215 | _T_5201; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24038.4]
  assign _T_5219 = _T_5217 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24040.4]
  assign _T_5220 = _T_5219 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24041.4]
  assign _T_5221 = _T_5206 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24046.4]
  assign _T_5222 = _T_5201 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24047.4]
  assign _T_5223 = _T_5221 | _T_5222; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24048.4]
  assign _T_5225 = _T_5223 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24050.4]
  assign _T_5226 = _T_5225 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24051.4]
  assign _T_5237 = _T_2494 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24068.4]
  assign _T_5238 = _T_2754 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24069.4]
  assign _T_5240 = _T_5238 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24071.4]
  assign _T_5242 = _T_5232 + _T_5237; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24073.4]
  assign _T_5243 = _T_5242 - _T_5240; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24074.4]
  assign _T_5244 = $unsigned(_T_5243); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24075.4]
  assign _T_5245 = _T_5244[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24076.4]
  assign _T_5246 = _T_5240 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24078.4]
  assign _T_5248 = _T_5246 | _T_5232; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24080.4]
  assign _T_5250 = _T_5248 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24082.4]
  assign _T_5251 = _T_5250 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24083.4]
  assign _T_5252 = _T_5237 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24088.4]
  assign _T_5253 = _T_5232 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24089.4]
  assign _T_5254 = _T_5252 | _T_5253; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24090.4]
  assign _T_5256 = _T_5254 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24092.4]
  assign _T_5257 = _T_5256 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24093.4]
  assign _T_5268 = _T_2495 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24110.4]
  assign _T_5269 = _T_2755 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24111.4]
  assign _T_5271 = _T_5269 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24113.4]
  assign _T_5273 = _T_5263 + _T_5268; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24115.4]
  assign _T_5274 = _T_5273 - _T_5271; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24116.4]
  assign _T_5275 = $unsigned(_T_5274); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24117.4]
  assign _T_5276 = _T_5275[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24118.4]
  assign _T_5277 = _T_5271 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24120.4]
  assign _T_5279 = _T_5277 | _T_5263; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24122.4]
  assign _T_5281 = _T_5279 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24124.4]
  assign _T_5282 = _T_5281 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24125.4]
  assign _T_5283 = _T_5268 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24130.4]
  assign _T_5284 = _T_5263 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24131.4]
  assign _T_5285 = _T_5283 | _T_5284; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24132.4]
  assign _T_5287 = _T_5285 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24134.4]
  assign _T_5288 = _T_5287 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24135.4]
  assign _T_5299 = _T_2496 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24152.4]
  assign _T_5300 = _T_2756 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24153.4]
  assign _T_5302 = _T_5300 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24155.4]
  assign _T_5304 = _T_5294 + _T_5299; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24157.4]
  assign _T_5305 = _T_5304 - _T_5302; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24158.4]
  assign _T_5306 = $unsigned(_T_5305); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24159.4]
  assign _T_5307 = _T_5306[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24160.4]
  assign _T_5308 = _T_5302 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24162.4]
  assign _T_5310 = _T_5308 | _T_5294; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24164.4]
  assign _T_5312 = _T_5310 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24166.4]
  assign _T_5313 = _T_5312 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24167.4]
  assign _T_5314 = _T_5299 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24172.4]
  assign _T_5315 = _T_5294 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24173.4]
  assign _T_5316 = _T_5314 | _T_5315; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24174.4]
  assign _T_5318 = _T_5316 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24176.4]
  assign _T_5319 = _T_5318 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24177.4]
  assign _T_5330 = _T_2497 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24194.4]
  assign _T_5331 = _T_2757 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24195.4]
  assign _T_5333 = _T_5331 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24197.4]
  assign _T_5335 = _T_5325 + _T_5330; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24199.4]
  assign _T_5336 = _T_5335 - _T_5333; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24200.4]
  assign _T_5337 = $unsigned(_T_5336); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24201.4]
  assign _T_5338 = _T_5337[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24202.4]
  assign _T_5339 = _T_5333 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24204.4]
  assign _T_5341 = _T_5339 | _T_5325; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24206.4]
  assign _T_5343 = _T_5341 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24208.4]
  assign _T_5344 = _T_5343 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24209.4]
  assign _T_5345 = _T_5330 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24214.4]
  assign _T_5346 = _T_5325 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24215.4]
  assign _T_5347 = _T_5345 | _T_5346; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24216.4]
  assign _T_5349 = _T_5347 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24218.4]
  assign _T_5350 = _T_5349 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24219.4]
  assign _T_5361 = _T_2498 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24236.4]
  assign _T_5362 = _T_2758 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24237.4]
  assign _T_5364 = _T_5362 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24239.4]
  assign _T_5366 = _T_5356 + _T_5361; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24241.4]
  assign _T_5367 = _T_5366 - _T_5364; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24242.4]
  assign _T_5368 = $unsigned(_T_5367); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24243.4]
  assign _T_5369 = _T_5368[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24244.4]
  assign _T_5370 = _T_5364 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24246.4]
  assign _T_5372 = _T_5370 | _T_5356; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24248.4]
  assign _T_5374 = _T_5372 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24250.4]
  assign _T_5375 = _T_5374 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24251.4]
  assign _T_5376 = _T_5361 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24256.4]
  assign _T_5377 = _T_5356 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24257.4]
  assign _T_5378 = _T_5376 | _T_5377; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24258.4]
  assign _T_5380 = _T_5378 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24260.4]
  assign _T_5381 = _T_5380 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24261.4]
  assign _T_5392 = _T_2499 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24278.4]
  assign _T_5393 = _T_2759 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24279.4]
  assign _T_5395 = _T_5393 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24281.4]
  assign _T_5397 = _T_5387 + _T_5392; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24283.4]
  assign _T_5398 = _T_5397 - _T_5395; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24284.4]
  assign _T_5399 = $unsigned(_T_5398); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24285.4]
  assign _T_5400 = _T_5399[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24286.4]
  assign _T_5401 = _T_5395 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24288.4]
  assign _T_5403 = _T_5401 | _T_5387; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24290.4]
  assign _T_5405 = _T_5403 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24292.4]
  assign _T_5406 = _T_5405 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24293.4]
  assign _T_5407 = _T_5392 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24298.4]
  assign _T_5408 = _T_5387 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24299.4]
  assign _T_5409 = _T_5407 | _T_5408; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24300.4]
  assign _T_5411 = _T_5409 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24302.4]
  assign _T_5412 = _T_5411 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24303.4]
  assign _T_5423 = _T_2500 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24320.4]
  assign _T_5424 = _T_2760 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24321.4]
  assign _T_5426 = _T_5424 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24323.4]
  assign _T_5428 = _T_5418 + _T_5423; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24325.4]
  assign _T_5429 = _T_5428 - _T_5426; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24326.4]
  assign _T_5430 = $unsigned(_T_5429); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24327.4]
  assign _T_5431 = _T_5430[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24328.4]
  assign _T_5432 = _T_5426 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24330.4]
  assign _T_5434 = _T_5432 | _T_5418; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24332.4]
  assign _T_5436 = _T_5434 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24334.4]
  assign _T_5437 = _T_5436 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24335.4]
  assign _T_5438 = _T_5423 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24340.4]
  assign _T_5439 = _T_5418 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24341.4]
  assign _T_5440 = _T_5438 | _T_5439; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24342.4]
  assign _T_5442 = _T_5440 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24344.4]
  assign _T_5443 = _T_5442 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24345.4]
  assign _T_5454 = _T_2501 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24362.4]
  assign _T_5455 = _T_2761 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24363.4]
  assign _T_5457 = _T_5455 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24365.4]
  assign _T_5459 = _T_5449 + _T_5454; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24367.4]
  assign _T_5460 = _T_5459 - _T_5457; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24368.4]
  assign _T_5461 = $unsigned(_T_5460); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24369.4]
  assign _T_5462 = _T_5461[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24370.4]
  assign _T_5463 = _T_5457 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24372.4]
  assign _T_5465 = _T_5463 | _T_5449; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24374.4]
  assign _T_5467 = _T_5465 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24376.4]
  assign _T_5468 = _T_5467 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24377.4]
  assign _T_5469 = _T_5454 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24382.4]
  assign _T_5470 = _T_5449 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24383.4]
  assign _T_5471 = _T_5469 | _T_5470; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24384.4]
  assign _T_5473 = _T_5471 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24386.4]
  assign _T_5474 = _T_5473 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24387.4]
  assign _T_5485 = _T_2502 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24404.4]
  assign _T_5486 = _T_2762 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24405.4]
  assign _T_5488 = _T_5486 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24407.4]
  assign _T_5490 = _T_5480 + _T_5485; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24409.4]
  assign _T_5491 = _T_5490 - _T_5488; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24410.4]
  assign _T_5492 = $unsigned(_T_5491); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24411.4]
  assign _T_5493 = _T_5492[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24412.4]
  assign _T_5494 = _T_5488 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24414.4]
  assign _T_5496 = _T_5494 | _T_5480; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24416.4]
  assign _T_5498 = _T_5496 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24418.4]
  assign _T_5499 = _T_5498 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24419.4]
  assign _T_5500 = _T_5485 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24424.4]
  assign _T_5501 = _T_5480 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24425.4]
  assign _T_5502 = _T_5500 | _T_5501; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24426.4]
  assign _T_5504 = _T_5502 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24428.4]
  assign _T_5505 = _T_5504 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24429.4]
  assign _T_5516 = _T_2503 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24446.4]
  assign _T_5517 = _T_2763 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24447.4]
  assign _T_5519 = _T_5517 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24449.4]
  assign _T_5521 = _T_5511 + _T_5516; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24451.4]
  assign _T_5522 = _T_5521 - _T_5519; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24452.4]
  assign _T_5523 = $unsigned(_T_5522); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24453.4]
  assign _T_5524 = _T_5523[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24454.4]
  assign _T_5525 = _T_5519 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24456.4]
  assign _T_5527 = _T_5525 | _T_5511; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24458.4]
  assign _T_5529 = _T_5527 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24460.4]
  assign _T_5530 = _T_5529 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24461.4]
  assign _T_5531 = _T_5516 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24466.4]
  assign _T_5532 = _T_5511 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24467.4]
  assign _T_5533 = _T_5531 | _T_5532; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24468.4]
  assign _T_5535 = _T_5533 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24470.4]
  assign _T_5536 = _T_5535 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24471.4]
  assign _T_5547 = _T_2504 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24488.4]
  assign _T_5548 = _T_2764 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24489.4]
  assign _T_5550 = _T_5548 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24491.4]
  assign _T_5552 = _T_5542 + _T_5547; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24493.4]
  assign _T_5553 = _T_5552 - _T_5550; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24494.4]
  assign _T_5554 = $unsigned(_T_5553); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24495.4]
  assign _T_5555 = _T_5554[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24496.4]
  assign _T_5556 = _T_5550 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24498.4]
  assign _T_5558 = _T_5556 | _T_5542; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24500.4]
  assign _T_5560 = _T_5558 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24502.4]
  assign _T_5561 = _T_5560 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24503.4]
  assign _T_5562 = _T_5547 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24508.4]
  assign _T_5563 = _T_5542 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24509.4]
  assign _T_5564 = _T_5562 | _T_5563; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24510.4]
  assign _T_5566 = _T_5564 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24512.4]
  assign _T_5567 = _T_5566 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24513.4]
  assign _T_5578 = _T_2505 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24530.4]
  assign _T_5579 = _T_2765 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24531.4]
  assign _T_5581 = _T_5579 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24533.4]
  assign _T_5583 = _T_5573 + _T_5578; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24535.4]
  assign _T_5584 = _T_5583 - _T_5581; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24536.4]
  assign _T_5585 = $unsigned(_T_5584); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24537.4]
  assign _T_5586 = _T_5585[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24538.4]
  assign _T_5587 = _T_5581 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24540.4]
  assign _T_5589 = _T_5587 | _T_5573; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24542.4]
  assign _T_5591 = _T_5589 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24544.4]
  assign _T_5592 = _T_5591 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24545.4]
  assign _T_5593 = _T_5578 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24550.4]
  assign _T_5594 = _T_5573 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24551.4]
  assign _T_5595 = _T_5593 | _T_5594; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24552.4]
  assign _T_5597 = _T_5595 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24554.4]
  assign _T_5598 = _T_5597 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24555.4]
  assign _T_5609 = _T_2506 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24572.4]
  assign _T_5610 = _T_2766 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24573.4]
  assign _T_5612 = _T_5610 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24575.4]
  assign _T_5614 = _T_5604 + _T_5609; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24577.4]
  assign _T_5615 = _T_5614 - _T_5612; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24578.4]
  assign _T_5616 = $unsigned(_T_5615); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24579.4]
  assign _T_5617 = _T_5616[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24580.4]
  assign _T_5618 = _T_5612 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24582.4]
  assign _T_5620 = _T_5618 | _T_5604; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24584.4]
  assign _T_5622 = _T_5620 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24586.4]
  assign _T_5623 = _T_5622 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24587.4]
  assign _T_5624 = _T_5609 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24592.4]
  assign _T_5625 = _T_5604 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24593.4]
  assign _T_5626 = _T_5624 | _T_5625; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24594.4]
  assign _T_5628 = _T_5626 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24596.4]
  assign _T_5629 = _T_5628 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24597.4]
  assign _T_5640 = _T_2507 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24614.4]
  assign _T_5641 = _T_2767 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24615.4]
  assign _T_5643 = _T_5641 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24617.4]
  assign _T_5645 = _T_5635 + _T_5640; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24619.4]
  assign _T_5646 = _T_5645 - _T_5643; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24620.4]
  assign _T_5647 = $unsigned(_T_5646); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24621.4]
  assign _T_5648 = _T_5647[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24622.4]
  assign _T_5649 = _T_5643 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24624.4]
  assign _T_5651 = _T_5649 | _T_5635; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24626.4]
  assign _T_5653 = _T_5651 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24628.4]
  assign _T_5654 = _T_5653 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24629.4]
  assign _T_5655 = _T_5640 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24634.4]
  assign _T_5656 = _T_5635 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24635.4]
  assign _T_5657 = _T_5655 | _T_5656; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24636.4]
  assign _T_5659 = _T_5657 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24638.4]
  assign _T_5660 = _T_5659 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24639.4]
  assign _T_5671 = _T_2508 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24656.4]
  assign _T_5672 = _T_2768 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24657.4]
  assign _T_5674 = _T_5672 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24659.4]
  assign _T_5676 = _T_5666 + _T_5671; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24661.4]
  assign _T_5677 = _T_5676 - _T_5674; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24662.4]
  assign _T_5678 = $unsigned(_T_5677); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24663.4]
  assign _T_5679 = _T_5678[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24664.4]
  assign _T_5680 = _T_5674 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24666.4]
  assign _T_5682 = _T_5680 | _T_5666; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24668.4]
  assign _T_5684 = _T_5682 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24670.4]
  assign _T_5685 = _T_5684 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24671.4]
  assign _T_5686 = _T_5671 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24676.4]
  assign _T_5687 = _T_5666 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24677.4]
  assign _T_5688 = _T_5686 | _T_5687; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24678.4]
  assign _T_5690 = _T_5688 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24680.4]
  assign _T_5691 = _T_5690 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24681.4]
  assign _T_5702 = _T_2509 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24698.4]
  assign _T_5703 = _T_2769 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24699.4]
  assign _T_5705 = _T_5703 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24701.4]
  assign _T_5707 = _T_5697 + _T_5702; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24703.4]
  assign _T_5708 = _T_5707 - _T_5705; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24704.4]
  assign _T_5709 = $unsigned(_T_5708); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24705.4]
  assign _T_5710 = _T_5709[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24706.4]
  assign _T_5711 = _T_5705 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24708.4]
  assign _T_5713 = _T_5711 | _T_5697; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24710.4]
  assign _T_5715 = _T_5713 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24712.4]
  assign _T_5716 = _T_5715 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24713.4]
  assign _T_5717 = _T_5702 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24718.4]
  assign _T_5718 = _T_5697 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24719.4]
  assign _T_5719 = _T_5717 | _T_5718; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24720.4]
  assign _T_5721 = _T_5719 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24722.4]
  assign _T_5722 = _T_5721 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24723.4]
  assign _T_5733 = _T_2510 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24740.4]
  assign _T_5734 = _T_2770 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24741.4]
  assign _T_5736 = _T_5734 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24743.4]
  assign _T_5738 = _T_5728 + _T_5733; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24745.4]
  assign _T_5739 = _T_5738 - _T_5736; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24746.4]
  assign _T_5740 = $unsigned(_T_5739); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24747.4]
  assign _T_5741 = _T_5740[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24748.4]
  assign _T_5742 = _T_5736 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24750.4]
  assign _T_5744 = _T_5742 | _T_5728; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24752.4]
  assign _T_5746 = _T_5744 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24754.4]
  assign _T_5747 = _T_5746 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24755.4]
  assign _T_5748 = _T_5733 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24760.4]
  assign _T_5749 = _T_5728 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24761.4]
  assign _T_5750 = _T_5748 | _T_5749; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24762.4]
  assign _T_5752 = _T_5750 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24764.4]
  assign _T_5753 = _T_5752 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24765.4]
  assign _T_5764 = _T_2511 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24782.4]
  assign _T_5765 = _T_2771 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24783.4]
  assign _T_5767 = _T_5765 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24785.4]
  assign _T_5769 = _T_5759 + _T_5764; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24787.4]
  assign _T_5770 = _T_5769 - _T_5767; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24788.4]
  assign _T_5771 = $unsigned(_T_5770); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24789.4]
  assign _T_5772 = _T_5771[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24790.4]
  assign _T_5773 = _T_5767 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24792.4]
  assign _T_5775 = _T_5773 | _T_5759; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24794.4]
  assign _T_5777 = _T_5775 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24796.4]
  assign _T_5778 = _T_5777 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24797.4]
  assign _T_5779 = _T_5764 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24802.4]
  assign _T_5780 = _T_5759 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24803.4]
  assign _T_5781 = _T_5779 | _T_5780; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24804.4]
  assign _T_5783 = _T_5781 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24806.4]
  assign _T_5784 = _T_5783 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24807.4]
  assign _T_5795 = _T_2512 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24824.4]
  assign _T_5796 = _T_2772 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24825.4]
  assign _T_5798 = _T_5796 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24827.4]
  assign _T_5800 = _T_5790 + _T_5795; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24829.4]
  assign _T_5801 = _T_5800 - _T_5798; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24830.4]
  assign _T_5802 = $unsigned(_T_5801); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24831.4]
  assign _T_5803 = _T_5802[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24832.4]
  assign _T_5804 = _T_5798 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24834.4]
  assign _T_5806 = _T_5804 | _T_5790; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24836.4]
  assign _T_5808 = _T_5806 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24838.4]
  assign _T_5809 = _T_5808 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24839.4]
  assign _T_5810 = _T_5795 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24844.4]
  assign _T_5811 = _T_5790 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24845.4]
  assign _T_5812 = _T_5810 | _T_5811; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24846.4]
  assign _T_5814 = _T_5812 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24848.4]
  assign _T_5815 = _T_5814 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24849.4]
  assign _T_5826 = _T_2513 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24866.4]
  assign _T_5827 = _T_2773 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24867.4]
  assign _T_5829 = _T_5827 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24869.4]
  assign _T_5831 = _T_5821 + _T_5826; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24871.4]
  assign _T_5832 = _T_5831 - _T_5829; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24872.4]
  assign _T_5833 = $unsigned(_T_5832); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24873.4]
  assign _T_5834 = _T_5833[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24874.4]
  assign _T_5835 = _T_5829 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24876.4]
  assign _T_5837 = _T_5835 | _T_5821; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24878.4]
  assign _T_5839 = _T_5837 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24880.4]
  assign _T_5840 = _T_5839 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24881.4]
  assign _T_5841 = _T_5826 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24886.4]
  assign _T_5842 = _T_5821 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24887.4]
  assign _T_5843 = _T_5841 | _T_5842; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24888.4]
  assign _T_5845 = _T_5843 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24890.4]
  assign _T_5846 = _T_5845 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24891.4]
  assign _T_5857 = _T_2514 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24908.4]
  assign _T_5858 = _T_2774 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24909.4]
  assign _T_5860 = _T_5858 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24911.4]
  assign _T_5862 = _T_5852 + _T_5857; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24913.4]
  assign _T_5863 = _T_5862 - _T_5860; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24914.4]
  assign _T_5864 = $unsigned(_T_5863); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24915.4]
  assign _T_5865 = _T_5864[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24916.4]
  assign _T_5866 = _T_5860 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24918.4]
  assign _T_5868 = _T_5866 | _T_5852; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24920.4]
  assign _T_5870 = _T_5868 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24922.4]
  assign _T_5871 = _T_5870 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24923.4]
  assign _T_5872 = _T_5857 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24928.4]
  assign _T_5873 = _T_5852 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24929.4]
  assign _T_5874 = _T_5872 | _T_5873; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24930.4]
  assign _T_5876 = _T_5874 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24932.4]
  assign _T_5877 = _T_5876 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24933.4]
  assign _T_5888 = _T_2515 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24950.4]
  assign _T_5889 = _T_2775 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24951.4]
  assign _T_5891 = _T_5889 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24953.4]
  assign _T_5893 = _T_5883 + _T_5888; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24955.4]
  assign _T_5894 = _T_5893 - _T_5891; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24956.4]
  assign _T_5895 = $unsigned(_T_5894); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24957.4]
  assign _T_5896 = _T_5895[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24958.4]
  assign _T_5897 = _T_5891 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@24960.4]
  assign _T_5899 = _T_5897 | _T_5883; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@24962.4]
  assign _T_5901 = _T_5899 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24964.4]
  assign _T_5902 = _T_5901 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24965.4]
  assign _T_5903 = _T_5888 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@24970.4]
  assign _T_5904 = _T_5883 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@24971.4]
  assign _T_5905 = _T_5903 | _T_5904; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@24972.4]
  assign _T_5907 = _T_5905 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24974.4]
  assign _T_5908 = _T_5907 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24975.4]
  assign _T_5919 = _T_2516 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@24992.4]
  assign _T_5920 = _T_2776 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@24993.4]
  assign _T_5922 = _T_5920 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@24995.4]
  assign _T_5924 = _T_5914 + _T_5919; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@24997.4]
  assign _T_5925 = _T_5924 - _T_5922; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24998.4]
  assign _T_5926 = $unsigned(_T_5925); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@24999.4]
  assign _T_5927 = _T_5926[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25000.4]
  assign _T_5928 = _T_5922 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25002.4]
  assign _T_5930 = _T_5928 | _T_5914; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25004.4]
  assign _T_5932 = _T_5930 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25006.4]
  assign _T_5933 = _T_5932 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25007.4]
  assign _T_5934 = _T_5919 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25012.4]
  assign _T_5935 = _T_5914 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25013.4]
  assign _T_5936 = _T_5934 | _T_5935; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25014.4]
  assign _T_5938 = _T_5936 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25016.4]
  assign _T_5939 = _T_5938 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25017.4]
  assign _T_5950 = _T_2517 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25034.4]
  assign _T_5951 = _T_2777 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25035.4]
  assign _T_5953 = _T_5951 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25037.4]
  assign _T_5955 = _T_5945 + _T_5950; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25039.4]
  assign _T_5956 = _T_5955 - _T_5953; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25040.4]
  assign _T_5957 = $unsigned(_T_5956); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25041.4]
  assign _T_5958 = _T_5957[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25042.4]
  assign _T_5959 = _T_5953 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25044.4]
  assign _T_5961 = _T_5959 | _T_5945; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25046.4]
  assign _T_5963 = _T_5961 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25048.4]
  assign _T_5964 = _T_5963 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25049.4]
  assign _T_5965 = _T_5950 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25054.4]
  assign _T_5966 = _T_5945 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25055.4]
  assign _T_5967 = _T_5965 | _T_5966; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25056.4]
  assign _T_5969 = _T_5967 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25058.4]
  assign _T_5970 = _T_5969 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25059.4]
  assign _T_5981 = _T_2518 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25076.4]
  assign _T_5982 = _T_2778 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25077.4]
  assign _T_5984 = _T_5982 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25079.4]
  assign _T_5986 = _T_5976 + _T_5981; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25081.4]
  assign _T_5987 = _T_5986 - _T_5984; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25082.4]
  assign _T_5988 = $unsigned(_T_5987); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25083.4]
  assign _T_5989 = _T_5988[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25084.4]
  assign _T_5990 = _T_5984 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25086.4]
  assign _T_5992 = _T_5990 | _T_5976; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25088.4]
  assign _T_5994 = _T_5992 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25090.4]
  assign _T_5995 = _T_5994 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25091.4]
  assign _T_5996 = _T_5981 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25096.4]
  assign _T_5997 = _T_5976 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25097.4]
  assign _T_5998 = _T_5996 | _T_5997; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25098.4]
  assign _T_6000 = _T_5998 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25100.4]
  assign _T_6001 = _T_6000 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25101.4]
  assign _T_6012 = _T_2519 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25118.4]
  assign _T_6013 = _T_2779 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25119.4]
  assign _T_6015 = _T_6013 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25121.4]
  assign _T_6017 = _T_6007 + _T_6012; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25123.4]
  assign _T_6018 = _T_6017 - _T_6015; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25124.4]
  assign _T_6019 = $unsigned(_T_6018); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25125.4]
  assign _T_6020 = _T_6019[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25126.4]
  assign _T_6021 = _T_6015 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25128.4]
  assign _T_6023 = _T_6021 | _T_6007; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25130.4]
  assign _T_6025 = _T_6023 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25132.4]
  assign _T_6026 = _T_6025 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25133.4]
  assign _T_6027 = _T_6012 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25138.4]
  assign _T_6028 = _T_6007 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25139.4]
  assign _T_6029 = _T_6027 | _T_6028; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25140.4]
  assign _T_6031 = _T_6029 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25142.4]
  assign _T_6032 = _T_6031 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25143.4]
  assign _T_6043 = _T_2520 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25160.4]
  assign _T_6044 = _T_2780 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25161.4]
  assign _T_6046 = _T_6044 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25163.4]
  assign _T_6048 = _T_6038 + _T_6043; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25165.4]
  assign _T_6049 = _T_6048 - _T_6046; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25166.4]
  assign _T_6050 = $unsigned(_T_6049); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25167.4]
  assign _T_6051 = _T_6050[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25168.4]
  assign _T_6052 = _T_6046 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25170.4]
  assign _T_6054 = _T_6052 | _T_6038; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25172.4]
  assign _T_6056 = _T_6054 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25174.4]
  assign _T_6057 = _T_6056 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25175.4]
  assign _T_6058 = _T_6043 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25180.4]
  assign _T_6059 = _T_6038 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25181.4]
  assign _T_6060 = _T_6058 | _T_6059; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25182.4]
  assign _T_6062 = _T_6060 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25184.4]
  assign _T_6063 = _T_6062 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25185.4]
  assign _T_6074 = _T_2521 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25202.4]
  assign _T_6075 = _T_2781 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25203.4]
  assign _T_6077 = _T_6075 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25205.4]
  assign _T_6079 = _T_6069 + _T_6074; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25207.4]
  assign _T_6080 = _T_6079 - _T_6077; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25208.4]
  assign _T_6081 = $unsigned(_T_6080); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25209.4]
  assign _T_6082 = _T_6081[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25210.4]
  assign _T_6083 = _T_6077 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25212.4]
  assign _T_6085 = _T_6083 | _T_6069; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25214.4]
  assign _T_6087 = _T_6085 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25216.4]
  assign _T_6088 = _T_6087 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25217.4]
  assign _T_6089 = _T_6074 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25222.4]
  assign _T_6090 = _T_6069 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25223.4]
  assign _T_6091 = _T_6089 | _T_6090; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25224.4]
  assign _T_6093 = _T_6091 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25226.4]
  assign _T_6094 = _T_6093 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25227.4]
  assign _T_6105 = _T_2522 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25244.4]
  assign _T_6106 = _T_2782 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25245.4]
  assign _T_6108 = _T_6106 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25247.4]
  assign _T_6110 = _T_6100 + _T_6105; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25249.4]
  assign _T_6111 = _T_6110 - _T_6108; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25250.4]
  assign _T_6112 = $unsigned(_T_6111); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25251.4]
  assign _T_6113 = _T_6112[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25252.4]
  assign _T_6114 = _T_6108 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25254.4]
  assign _T_6116 = _T_6114 | _T_6100; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25256.4]
  assign _T_6118 = _T_6116 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25258.4]
  assign _T_6119 = _T_6118 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25259.4]
  assign _T_6120 = _T_6105 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25264.4]
  assign _T_6121 = _T_6100 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25265.4]
  assign _T_6122 = _T_6120 | _T_6121; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25266.4]
  assign _T_6124 = _T_6122 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25268.4]
  assign _T_6125 = _T_6124 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25269.4]
  assign _T_6136 = _T_2523 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25286.4]
  assign _T_6137 = _T_2783 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25287.4]
  assign _T_6139 = _T_6137 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25289.4]
  assign _T_6141 = _T_6131 + _T_6136; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25291.4]
  assign _T_6142 = _T_6141 - _T_6139; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25292.4]
  assign _T_6143 = $unsigned(_T_6142); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25293.4]
  assign _T_6144 = _T_6143[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25294.4]
  assign _T_6145 = _T_6139 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25296.4]
  assign _T_6147 = _T_6145 | _T_6131; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25298.4]
  assign _T_6149 = _T_6147 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25300.4]
  assign _T_6150 = _T_6149 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25301.4]
  assign _T_6151 = _T_6136 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25306.4]
  assign _T_6152 = _T_6131 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25307.4]
  assign _T_6153 = _T_6151 | _T_6152; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25308.4]
  assign _T_6155 = _T_6153 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25310.4]
  assign _T_6156 = _T_6155 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25311.4]
  assign _T_6167 = _T_2524 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25328.4]
  assign _T_6168 = _T_2784 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25329.4]
  assign _T_6170 = _T_6168 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25331.4]
  assign _T_6172 = _T_6162 + _T_6167; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25333.4]
  assign _T_6173 = _T_6172 - _T_6170; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25334.4]
  assign _T_6174 = $unsigned(_T_6173); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25335.4]
  assign _T_6175 = _T_6174[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25336.4]
  assign _T_6176 = _T_6170 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25338.4]
  assign _T_6178 = _T_6176 | _T_6162; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25340.4]
  assign _T_6180 = _T_6178 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25342.4]
  assign _T_6181 = _T_6180 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25343.4]
  assign _T_6182 = _T_6167 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25348.4]
  assign _T_6183 = _T_6162 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25349.4]
  assign _T_6184 = _T_6182 | _T_6183; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25350.4]
  assign _T_6186 = _T_6184 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25352.4]
  assign _T_6187 = _T_6186 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25353.4]
  assign _T_6198 = _T_2525 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25370.4]
  assign _T_6199 = _T_2785 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25371.4]
  assign _T_6201 = _T_6199 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25373.4]
  assign _T_6203 = _T_6193 + _T_6198; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25375.4]
  assign _T_6204 = _T_6203 - _T_6201; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25376.4]
  assign _T_6205 = $unsigned(_T_6204); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25377.4]
  assign _T_6206 = _T_6205[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25378.4]
  assign _T_6207 = _T_6201 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25380.4]
  assign _T_6209 = _T_6207 | _T_6193; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25382.4]
  assign _T_6211 = _T_6209 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25384.4]
  assign _T_6212 = _T_6211 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25385.4]
  assign _T_6213 = _T_6198 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25390.4]
  assign _T_6214 = _T_6193 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25391.4]
  assign _T_6215 = _T_6213 | _T_6214; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25392.4]
  assign _T_6217 = _T_6215 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25394.4]
  assign _T_6218 = _T_6217 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25395.4]
  assign _T_6229 = _T_2526 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25412.4]
  assign _T_6230 = _T_2786 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25413.4]
  assign _T_6232 = _T_6230 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25415.4]
  assign _T_6234 = _T_6224 + _T_6229; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25417.4]
  assign _T_6235 = _T_6234 - _T_6232; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25418.4]
  assign _T_6236 = $unsigned(_T_6235); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25419.4]
  assign _T_6237 = _T_6236[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25420.4]
  assign _T_6238 = _T_6232 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25422.4]
  assign _T_6240 = _T_6238 | _T_6224; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25424.4]
  assign _T_6242 = _T_6240 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25426.4]
  assign _T_6243 = _T_6242 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25427.4]
  assign _T_6244 = _T_6229 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25432.4]
  assign _T_6245 = _T_6224 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25433.4]
  assign _T_6246 = _T_6244 | _T_6245; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25434.4]
  assign _T_6248 = _T_6246 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25436.4]
  assign _T_6249 = _T_6248 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25437.4]
  assign _T_6260 = _T_2527 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25454.4]
  assign _T_6261 = _T_2787 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25455.4]
  assign _T_6263 = _T_6261 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25457.4]
  assign _T_6265 = _T_6255 + _T_6260; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25459.4]
  assign _T_6266 = _T_6265 - _T_6263; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25460.4]
  assign _T_6267 = $unsigned(_T_6266); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25461.4]
  assign _T_6268 = _T_6267[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25462.4]
  assign _T_6269 = _T_6263 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25464.4]
  assign _T_6271 = _T_6269 | _T_6255; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25466.4]
  assign _T_6273 = _T_6271 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25468.4]
  assign _T_6274 = _T_6273 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25469.4]
  assign _T_6275 = _T_6260 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25474.4]
  assign _T_6276 = _T_6255 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25475.4]
  assign _T_6277 = _T_6275 | _T_6276; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25476.4]
  assign _T_6279 = _T_6277 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25478.4]
  assign _T_6280 = _T_6279 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25479.4]
  assign _T_6291 = _T_2528 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25496.4]
  assign _T_6292 = _T_2788 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25497.4]
  assign _T_6294 = _T_6292 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25499.4]
  assign _T_6296 = _T_6286 + _T_6291; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25501.4]
  assign _T_6297 = _T_6296 - _T_6294; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25502.4]
  assign _T_6298 = $unsigned(_T_6297); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25503.4]
  assign _T_6299 = _T_6298[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25504.4]
  assign _T_6300 = _T_6294 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25506.4]
  assign _T_6302 = _T_6300 | _T_6286; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25508.4]
  assign _T_6304 = _T_6302 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25510.4]
  assign _T_6305 = _T_6304 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25511.4]
  assign _T_6306 = _T_6291 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25516.4]
  assign _T_6307 = _T_6286 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25517.4]
  assign _T_6308 = _T_6306 | _T_6307; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25518.4]
  assign _T_6310 = _T_6308 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25520.4]
  assign _T_6311 = _T_6310 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25521.4]
  assign _T_6322 = _T_2529 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25538.4]
  assign _T_6323 = _T_2789 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25539.4]
  assign _T_6325 = _T_6323 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25541.4]
  assign _T_6327 = _T_6317 + _T_6322; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25543.4]
  assign _T_6328 = _T_6327 - _T_6325; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25544.4]
  assign _T_6329 = $unsigned(_T_6328); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25545.4]
  assign _T_6330 = _T_6329[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25546.4]
  assign _T_6331 = _T_6325 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25548.4]
  assign _T_6333 = _T_6331 | _T_6317; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25550.4]
  assign _T_6335 = _T_6333 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25552.4]
  assign _T_6336 = _T_6335 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25553.4]
  assign _T_6337 = _T_6322 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25558.4]
  assign _T_6338 = _T_6317 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25559.4]
  assign _T_6339 = _T_6337 | _T_6338; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25560.4]
  assign _T_6341 = _T_6339 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25562.4]
  assign _T_6342 = _T_6341 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25563.4]
  assign _T_6353 = _T_2530 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25580.4]
  assign _T_6354 = _T_2790 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25581.4]
  assign _T_6356 = _T_6354 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25583.4]
  assign _T_6358 = _T_6348 + _T_6353; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25585.4]
  assign _T_6359 = _T_6358 - _T_6356; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25586.4]
  assign _T_6360 = $unsigned(_T_6359); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25587.4]
  assign _T_6361 = _T_6360[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25588.4]
  assign _T_6362 = _T_6356 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25590.4]
  assign _T_6364 = _T_6362 | _T_6348; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25592.4]
  assign _T_6366 = _T_6364 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25594.4]
  assign _T_6367 = _T_6366 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25595.4]
  assign _T_6368 = _T_6353 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25600.4]
  assign _T_6369 = _T_6348 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25601.4]
  assign _T_6370 = _T_6368 | _T_6369; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25602.4]
  assign _T_6372 = _T_6370 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25604.4]
  assign _T_6373 = _T_6372 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25605.4]
  assign _T_6384 = _T_2531 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25622.4]
  assign _T_6385 = _T_2791 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25623.4]
  assign _T_6387 = _T_6385 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25625.4]
  assign _T_6389 = _T_6379 + _T_6384; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25627.4]
  assign _T_6390 = _T_6389 - _T_6387; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25628.4]
  assign _T_6391 = $unsigned(_T_6390); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25629.4]
  assign _T_6392 = _T_6391[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25630.4]
  assign _T_6393 = _T_6387 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25632.4]
  assign _T_6395 = _T_6393 | _T_6379; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25634.4]
  assign _T_6397 = _T_6395 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25636.4]
  assign _T_6398 = _T_6397 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25637.4]
  assign _T_6399 = _T_6384 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25642.4]
  assign _T_6400 = _T_6379 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25643.4]
  assign _T_6401 = _T_6399 | _T_6400; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25644.4]
  assign _T_6403 = _T_6401 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25646.4]
  assign _T_6404 = _T_6403 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25647.4]
  assign _T_6415 = _T_2532 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25664.4]
  assign _T_6416 = _T_2792 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25665.4]
  assign _T_6418 = _T_6416 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25667.4]
  assign _T_6420 = _T_6410 + _T_6415; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25669.4]
  assign _T_6421 = _T_6420 - _T_6418; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25670.4]
  assign _T_6422 = $unsigned(_T_6421); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25671.4]
  assign _T_6423 = _T_6422[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25672.4]
  assign _T_6424 = _T_6418 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25674.4]
  assign _T_6426 = _T_6424 | _T_6410; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25676.4]
  assign _T_6428 = _T_6426 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25678.4]
  assign _T_6429 = _T_6428 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25679.4]
  assign _T_6430 = _T_6415 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25684.4]
  assign _T_6431 = _T_6410 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25685.4]
  assign _T_6432 = _T_6430 | _T_6431; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25686.4]
  assign _T_6434 = _T_6432 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25688.4]
  assign _T_6435 = _T_6434 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25689.4]
  assign _T_6446 = _T_2533 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25706.4]
  assign _T_6447 = _T_2793 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25707.4]
  assign _T_6449 = _T_6447 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25709.4]
  assign _T_6451 = _T_6441 + _T_6446; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25711.4]
  assign _T_6452 = _T_6451 - _T_6449; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25712.4]
  assign _T_6453 = $unsigned(_T_6452); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25713.4]
  assign _T_6454 = _T_6453[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25714.4]
  assign _T_6455 = _T_6449 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25716.4]
  assign _T_6457 = _T_6455 | _T_6441; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25718.4]
  assign _T_6459 = _T_6457 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25720.4]
  assign _T_6460 = _T_6459 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25721.4]
  assign _T_6461 = _T_6446 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25726.4]
  assign _T_6462 = _T_6441 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25727.4]
  assign _T_6463 = _T_6461 | _T_6462; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25728.4]
  assign _T_6465 = _T_6463 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25730.4]
  assign _T_6466 = _T_6465 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25731.4]
  assign _T_6477 = _T_2534 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25748.4]
  assign _T_6478 = _T_2794 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25749.4]
  assign _T_6480 = _T_6478 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25751.4]
  assign _T_6482 = _T_6472 + _T_6477; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25753.4]
  assign _T_6483 = _T_6482 - _T_6480; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25754.4]
  assign _T_6484 = $unsigned(_T_6483); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25755.4]
  assign _T_6485 = _T_6484[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25756.4]
  assign _T_6486 = _T_6480 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25758.4]
  assign _T_6488 = _T_6486 | _T_6472; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25760.4]
  assign _T_6490 = _T_6488 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25762.4]
  assign _T_6491 = _T_6490 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25763.4]
  assign _T_6492 = _T_6477 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25768.4]
  assign _T_6493 = _T_6472 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25769.4]
  assign _T_6494 = _T_6492 | _T_6493; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25770.4]
  assign _T_6496 = _T_6494 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25772.4]
  assign _T_6497 = _T_6496 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25773.4]
  assign _T_6508 = _T_2535 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25790.4]
  assign _T_6509 = _T_2795 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25791.4]
  assign _T_6511 = _T_6509 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25793.4]
  assign _T_6513 = _T_6503 + _T_6508; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25795.4]
  assign _T_6514 = _T_6513 - _T_6511; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25796.4]
  assign _T_6515 = $unsigned(_T_6514); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25797.4]
  assign _T_6516 = _T_6515[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25798.4]
  assign _T_6517 = _T_6511 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25800.4]
  assign _T_6519 = _T_6517 | _T_6503; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25802.4]
  assign _T_6521 = _T_6519 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25804.4]
  assign _T_6522 = _T_6521 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25805.4]
  assign _T_6523 = _T_6508 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25810.4]
  assign _T_6524 = _T_6503 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25811.4]
  assign _T_6525 = _T_6523 | _T_6524; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25812.4]
  assign _T_6527 = _T_6525 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25814.4]
  assign _T_6528 = _T_6527 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25815.4]
  assign _T_6539 = _T_2536 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25832.4]
  assign _T_6540 = _T_2796 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25833.4]
  assign _T_6542 = _T_6540 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25835.4]
  assign _T_6544 = _T_6534 + _T_6539; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25837.4]
  assign _T_6545 = _T_6544 - _T_6542; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25838.4]
  assign _T_6546 = $unsigned(_T_6545); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25839.4]
  assign _T_6547 = _T_6546[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25840.4]
  assign _T_6548 = _T_6542 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25842.4]
  assign _T_6550 = _T_6548 | _T_6534; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25844.4]
  assign _T_6552 = _T_6550 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25846.4]
  assign _T_6553 = _T_6552 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25847.4]
  assign _T_6554 = _T_6539 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25852.4]
  assign _T_6555 = _T_6534 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25853.4]
  assign _T_6556 = _T_6554 | _T_6555; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25854.4]
  assign _T_6558 = _T_6556 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25856.4]
  assign _T_6559 = _T_6558 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25857.4]
  assign _T_6570 = _T_2537 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25874.4]
  assign _T_6571 = _T_2797 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25875.4]
  assign _T_6573 = _T_6571 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25877.4]
  assign _T_6575 = _T_6565 + _T_6570; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25879.4]
  assign _T_6576 = _T_6575 - _T_6573; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25880.4]
  assign _T_6577 = $unsigned(_T_6576); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25881.4]
  assign _T_6578 = _T_6577[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25882.4]
  assign _T_6579 = _T_6573 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25884.4]
  assign _T_6581 = _T_6579 | _T_6565; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25886.4]
  assign _T_6583 = _T_6581 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25888.4]
  assign _T_6584 = _T_6583 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25889.4]
  assign _T_6585 = _T_6570 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25894.4]
  assign _T_6586 = _T_6565 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25895.4]
  assign _T_6587 = _T_6585 | _T_6586; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25896.4]
  assign _T_6589 = _T_6587 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25898.4]
  assign _T_6590 = _T_6589 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25899.4]
  assign _T_6601 = _T_2538 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25916.4]
  assign _T_6602 = _T_2798 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25917.4]
  assign _T_6604 = _T_6602 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25919.4]
  assign _T_6606 = _T_6596 + _T_6601; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25921.4]
  assign _T_6607 = _T_6606 - _T_6604; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25922.4]
  assign _T_6608 = $unsigned(_T_6607); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25923.4]
  assign _T_6609 = _T_6608[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25924.4]
  assign _T_6610 = _T_6604 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25926.4]
  assign _T_6612 = _T_6610 | _T_6596; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25928.4]
  assign _T_6614 = _T_6612 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25930.4]
  assign _T_6615 = _T_6614 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25931.4]
  assign _T_6616 = _T_6601 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25936.4]
  assign _T_6617 = _T_6596 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25937.4]
  assign _T_6618 = _T_6616 | _T_6617; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25938.4]
  assign _T_6620 = _T_6618 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25940.4]
  assign _T_6621 = _T_6620 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25941.4]
  assign _T_6632 = _T_2539 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@25958.4]
  assign _T_6633 = _T_2799 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@25959.4]
  assign _T_6635 = _T_6633 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@25961.4]
  assign _T_6637 = _T_6627 + _T_6632; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@25963.4]
  assign _T_6638 = _T_6637 - _T_6635; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25964.4]
  assign _T_6639 = $unsigned(_T_6638); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25965.4]
  assign _T_6640 = _T_6639[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@25966.4]
  assign _T_6641 = _T_6635 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@25968.4]
  assign _T_6643 = _T_6641 | _T_6627; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@25970.4]
  assign _T_6645 = _T_6643 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25972.4]
  assign _T_6646 = _T_6645 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25973.4]
  assign _T_6647 = _T_6632 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@25978.4]
  assign _T_6648 = _T_6627 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@25979.4]
  assign _T_6649 = _T_6647 | _T_6648; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@25980.4]
  assign _T_6651 = _T_6649 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25982.4]
  assign _T_6652 = _T_6651 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25983.4]
  assign _T_6663 = _T_2540 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26000.4]
  assign _T_6664 = _T_2800 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26001.4]
  assign _T_6666 = _T_6664 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26003.4]
  assign _T_6668 = _T_6658 + _T_6663; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26005.4]
  assign _T_6669 = _T_6668 - _T_6666; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26006.4]
  assign _T_6670 = $unsigned(_T_6669); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26007.4]
  assign _T_6671 = _T_6670[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26008.4]
  assign _T_6672 = _T_6666 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26010.4]
  assign _T_6674 = _T_6672 | _T_6658; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26012.4]
  assign _T_6676 = _T_6674 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26014.4]
  assign _T_6677 = _T_6676 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26015.4]
  assign _T_6678 = _T_6663 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26020.4]
  assign _T_6679 = _T_6658 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26021.4]
  assign _T_6680 = _T_6678 | _T_6679; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26022.4]
  assign _T_6682 = _T_6680 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26024.4]
  assign _T_6683 = _T_6682 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26025.4]
  assign _T_6694 = _T_2541 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26042.4]
  assign _T_6695 = _T_2801 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26043.4]
  assign _T_6697 = _T_6695 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26045.4]
  assign _T_6699 = _T_6689 + _T_6694; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26047.4]
  assign _T_6700 = _T_6699 - _T_6697; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26048.4]
  assign _T_6701 = $unsigned(_T_6700); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26049.4]
  assign _T_6702 = _T_6701[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26050.4]
  assign _T_6703 = _T_6697 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26052.4]
  assign _T_6705 = _T_6703 | _T_6689; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26054.4]
  assign _T_6707 = _T_6705 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26056.4]
  assign _T_6708 = _T_6707 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26057.4]
  assign _T_6709 = _T_6694 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26062.4]
  assign _T_6710 = _T_6689 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26063.4]
  assign _T_6711 = _T_6709 | _T_6710; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26064.4]
  assign _T_6713 = _T_6711 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26066.4]
  assign _T_6714 = _T_6713 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26067.4]
  assign _T_6725 = _T_2542 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26084.4]
  assign _T_6726 = _T_2802 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26085.4]
  assign _T_6728 = _T_6726 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26087.4]
  assign _T_6730 = _T_6720 + _T_6725; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26089.4]
  assign _T_6731 = _T_6730 - _T_6728; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26090.4]
  assign _T_6732 = $unsigned(_T_6731); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26091.4]
  assign _T_6733 = _T_6732[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26092.4]
  assign _T_6734 = _T_6728 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26094.4]
  assign _T_6736 = _T_6734 | _T_6720; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26096.4]
  assign _T_6738 = _T_6736 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26098.4]
  assign _T_6739 = _T_6738 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26099.4]
  assign _T_6740 = _T_6725 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26104.4]
  assign _T_6741 = _T_6720 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26105.4]
  assign _T_6742 = _T_6740 | _T_6741; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26106.4]
  assign _T_6744 = _T_6742 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26108.4]
  assign _T_6745 = _T_6744 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26109.4]
  assign _T_6756 = _T_2543 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26126.4]
  assign _T_6757 = _T_2803 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26127.4]
  assign _T_6759 = _T_6757 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26129.4]
  assign _T_6761 = _T_6751 + _T_6756; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26131.4]
  assign _T_6762 = _T_6761 - _T_6759; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26132.4]
  assign _T_6763 = $unsigned(_T_6762); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26133.4]
  assign _T_6764 = _T_6763[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26134.4]
  assign _T_6765 = _T_6759 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26136.4]
  assign _T_6767 = _T_6765 | _T_6751; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26138.4]
  assign _T_6769 = _T_6767 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26140.4]
  assign _T_6770 = _T_6769 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26141.4]
  assign _T_6771 = _T_6756 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26146.4]
  assign _T_6772 = _T_6751 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26147.4]
  assign _T_6773 = _T_6771 | _T_6772; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26148.4]
  assign _T_6775 = _T_6773 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26150.4]
  assign _T_6776 = _T_6775 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26151.4]
  assign _T_6787 = _T_2544 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26168.4]
  assign _T_6788 = _T_2804 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26169.4]
  assign _T_6790 = _T_6788 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26171.4]
  assign _T_6792 = _T_6782 + _T_6787; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26173.4]
  assign _T_6793 = _T_6792 - _T_6790; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26174.4]
  assign _T_6794 = $unsigned(_T_6793); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26175.4]
  assign _T_6795 = _T_6794[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26176.4]
  assign _T_6796 = _T_6790 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26178.4]
  assign _T_6798 = _T_6796 | _T_6782; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26180.4]
  assign _T_6800 = _T_6798 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26182.4]
  assign _T_6801 = _T_6800 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26183.4]
  assign _T_6802 = _T_6787 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26188.4]
  assign _T_6803 = _T_6782 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26189.4]
  assign _T_6804 = _T_6802 | _T_6803; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26190.4]
  assign _T_6806 = _T_6804 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26192.4]
  assign _T_6807 = _T_6806 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26193.4]
  assign _T_6818 = _T_2545 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26210.4]
  assign _T_6819 = _T_2805 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26211.4]
  assign _T_6821 = _T_6819 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26213.4]
  assign _T_6823 = _T_6813 + _T_6818; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26215.4]
  assign _T_6824 = _T_6823 - _T_6821; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26216.4]
  assign _T_6825 = $unsigned(_T_6824); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26217.4]
  assign _T_6826 = _T_6825[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26218.4]
  assign _T_6827 = _T_6821 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26220.4]
  assign _T_6829 = _T_6827 | _T_6813; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26222.4]
  assign _T_6831 = _T_6829 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26224.4]
  assign _T_6832 = _T_6831 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26225.4]
  assign _T_6833 = _T_6818 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26230.4]
  assign _T_6834 = _T_6813 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26231.4]
  assign _T_6835 = _T_6833 | _T_6834; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26232.4]
  assign _T_6837 = _T_6835 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26234.4]
  assign _T_6838 = _T_6837 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26235.4]
  assign _T_6849 = _T_2546 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26252.4]
  assign _T_6850 = _T_2806 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26253.4]
  assign _T_6852 = _T_6850 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26255.4]
  assign _T_6854 = _T_6844 + _T_6849; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26257.4]
  assign _T_6855 = _T_6854 - _T_6852; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26258.4]
  assign _T_6856 = $unsigned(_T_6855); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26259.4]
  assign _T_6857 = _T_6856[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26260.4]
  assign _T_6858 = _T_6852 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26262.4]
  assign _T_6860 = _T_6858 | _T_6844; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26264.4]
  assign _T_6862 = _T_6860 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26266.4]
  assign _T_6863 = _T_6862 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26267.4]
  assign _T_6864 = _T_6849 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26272.4]
  assign _T_6865 = _T_6844 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26273.4]
  assign _T_6866 = _T_6864 | _T_6865; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26274.4]
  assign _T_6868 = _T_6866 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26276.4]
  assign _T_6869 = _T_6868 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26277.4]
  assign _T_6880 = _T_2547 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26294.4]
  assign _T_6881 = _T_2807 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26295.4]
  assign _T_6883 = _T_6881 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26297.4]
  assign _T_6885 = _T_6875 + _T_6880; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26299.4]
  assign _T_6886 = _T_6885 - _T_6883; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26300.4]
  assign _T_6887 = $unsigned(_T_6886); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26301.4]
  assign _T_6888 = _T_6887[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26302.4]
  assign _T_6889 = _T_6883 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26304.4]
  assign _T_6891 = _T_6889 | _T_6875; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26306.4]
  assign _T_6893 = _T_6891 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26308.4]
  assign _T_6894 = _T_6893 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26309.4]
  assign _T_6895 = _T_6880 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26314.4]
  assign _T_6896 = _T_6875 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26315.4]
  assign _T_6897 = _T_6895 | _T_6896; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26316.4]
  assign _T_6899 = _T_6897 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26318.4]
  assign _T_6900 = _T_6899 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26319.4]
  assign _T_6911 = _T_2548 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26336.4]
  assign _T_6912 = _T_2808 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26337.4]
  assign _T_6914 = _T_6912 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26339.4]
  assign _T_6916 = _T_6906 + _T_6911; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26341.4]
  assign _T_6917 = _T_6916 - _T_6914; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26342.4]
  assign _T_6918 = $unsigned(_T_6917); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26343.4]
  assign _T_6919 = _T_6918[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26344.4]
  assign _T_6920 = _T_6914 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26346.4]
  assign _T_6922 = _T_6920 | _T_6906; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26348.4]
  assign _T_6924 = _T_6922 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26350.4]
  assign _T_6925 = _T_6924 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26351.4]
  assign _T_6926 = _T_6911 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26356.4]
  assign _T_6927 = _T_6906 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26357.4]
  assign _T_6928 = _T_6926 | _T_6927; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26358.4]
  assign _T_6930 = _T_6928 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26360.4]
  assign _T_6931 = _T_6930 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26361.4]
  assign _T_6942 = _T_2549 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26378.4]
  assign _T_6943 = _T_2809 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26379.4]
  assign _T_6945 = _T_6943 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26381.4]
  assign _T_6947 = _T_6937 + _T_6942; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26383.4]
  assign _T_6948 = _T_6947 - _T_6945; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26384.4]
  assign _T_6949 = $unsigned(_T_6948); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26385.4]
  assign _T_6950 = _T_6949[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26386.4]
  assign _T_6951 = _T_6945 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26388.4]
  assign _T_6953 = _T_6951 | _T_6937; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26390.4]
  assign _T_6955 = _T_6953 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26392.4]
  assign _T_6956 = _T_6955 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26393.4]
  assign _T_6957 = _T_6942 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26398.4]
  assign _T_6958 = _T_6937 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26399.4]
  assign _T_6959 = _T_6957 | _T_6958; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26400.4]
  assign _T_6961 = _T_6959 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26402.4]
  assign _T_6962 = _T_6961 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26403.4]
  assign _T_6973 = _T_2550 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26420.4]
  assign _T_6974 = _T_2810 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26421.4]
  assign _T_6976 = _T_6974 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26423.4]
  assign _T_6978 = _T_6968 + _T_6973; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26425.4]
  assign _T_6979 = _T_6978 - _T_6976; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26426.4]
  assign _T_6980 = $unsigned(_T_6979); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26427.4]
  assign _T_6981 = _T_6980[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26428.4]
  assign _T_6982 = _T_6976 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26430.4]
  assign _T_6984 = _T_6982 | _T_6968; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26432.4]
  assign _T_6986 = _T_6984 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26434.4]
  assign _T_6987 = _T_6986 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26435.4]
  assign _T_6988 = _T_6973 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26440.4]
  assign _T_6989 = _T_6968 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26441.4]
  assign _T_6990 = _T_6988 | _T_6989; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26442.4]
  assign _T_6992 = _T_6990 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26444.4]
  assign _T_6993 = _T_6992 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26445.4]
  assign _T_7004 = _T_2551 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26462.4]
  assign _T_7005 = _T_2811 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26463.4]
  assign _T_7007 = _T_7005 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26465.4]
  assign _T_7009 = _T_6999 + _T_7004; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26467.4]
  assign _T_7010 = _T_7009 - _T_7007; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26468.4]
  assign _T_7011 = $unsigned(_T_7010); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26469.4]
  assign _T_7012 = _T_7011[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26470.4]
  assign _T_7013 = _T_7007 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26472.4]
  assign _T_7015 = _T_7013 | _T_6999; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26474.4]
  assign _T_7017 = _T_7015 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26476.4]
  assign _T_7018 = _T_7017 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26477.4]
  assign _T_7019 = _T_7004 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26482.4]
  assign _T_7020 = _T_6999 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26483.4]
  assign _T_7021 = _T_7019 | _T_7020; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26484.4]
  assign _T_7023 = _T_7021 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26486.4]
  assign _T_7024 = _T_7023 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26487.4]
  assign _T_7035 = _T_2552 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26504.4]
  assign _T_7036 = _T_2812 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26505.4]
  assign _T_7038 = _T_7036 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26507.4]
  assign _T_7040 = _T_7030 + _T_7035; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26509.4]
  assign _T_7041 = _T_7040 - _T_7038; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26510.4]
  assign _T_7042 = $unsigned(_T_7041); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26511.4]
  assign _T_7043 = _T_7042[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26512.4]
  assign _T_7044 = _T_7038 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26514.4]
  assign _T_7046 = _T_7044 | _T_7030; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26516.4]
  assign _T_7048 = _T_7046 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26518.4]
  assign _T_7049 = _T_7048 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26519.4]
  assign _T_7050 = _T_7035 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26524.4]
  assign _T_7051 = _T_7030 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26525.4]
  assign _T_7052 = _T_7050 | _T_7051; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26526.4]
  assign _T_7054 = _T_7052 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26528.4]
  assign _T_7055 = _T_7054 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26529.4]
  assign _T_7066 = _T_2553 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26546.4]
  assign _T_7067 = _T_2813 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26547.4]
  assign _T_7069 = _T_7067 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26549.4]
  assign _T_7071 = _T_7061 + _T_7066; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26551.4]
  assign _T_7072 = _T_7071 - _T_7069; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26552.4]
  assign _T_7073 = $unsigned(_T_7072); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26553.4]
  assign _T_7074 = _T_7073[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26554.4]
  assign _T_7075 = _T_7069 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26556.4]
  assign _T_7077 = _T_7075 | _T_7061; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26558.4]
  assign _T_7079 = _T_7077 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26560.4]
  assign _T_7080 = _T_7079 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26561.4]
  assign _T_7081 = _T_7066 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26566.4]
  assign _T_7082 = _T_7061 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26567.4]
  assign _T_7083 = _T_7081 | _T_7082; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26568.4]
  assign _T_7085 = _T_7083 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26570.4]
  assign _T_7086 = _T_7085 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26571.4]
  assign _T_7097 = _T_2554 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26588.4]
  assign _T_7098 = _T_2814 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26589.4]
  assign _T_7100 = _T_7098 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26591.4]
  assign _T_7102 = _T_7092 + _T_7097; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26593.4]
  assign _T_7103 = _T_7102 - _T_7100; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26594.4]
  assign _T_7104 = $unsigned(_T_7103); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26595.4]
  assign _T_7105 = _T_7104[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26596.4]
  assign _T_7106 = _T_7100 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26598.4]
  assign _T_7108 = _T_7106 | _T_7092; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26600.4]
  assign _T_7110 = _T_7108 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26602.4]
  assign _T_7111 = _T_7110 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26603.4]
  assign _T_7112 = _T_7097 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26608.4]
  assign _T_7113 = _T_7092 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26609.4]
  assign _T_7114 = _T_7112 | _T_7113; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26610.4]
  assign _T_7116 = _T_7114 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26612.4]
  assign _T_7117 = _T_7116 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26613.4]
  assign _T_7128 = _T_2555 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26630.4]
  assign _T_7129 = _T_2815 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26631.4]
  assign _T_7131 = _T_7129 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26633.4]
  assign _T_7133 = _T_7123 + _T_7128; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26635.4]
  assign _T_7134 = _T_7133 - _T_7131; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26636.4]
  assign _T_7135 = $unsigned(_T_7134); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26637.4]
  assign _T_7136 = _T_7135[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26638.4]
  assign _T_7137 = _T_7131 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26640.4]
  assign _T_7139 = _T_7137 | _T_7123; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26642.4]
  assign _T_7141 = _T_7139 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26644.4]
  assign _T_7142 = _T_7141 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26645.4]
  assign _T_7143 = _T_7128 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26650.4]
  assign _T_7144 = _T_7123 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26651.4]
  assign _T_7145 = _T_7143 | _T_7144; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26652.4]
  assign _T_7147 = _T_7145 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26654.4]
  assign _T_7148 = _T_7147 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26655.4]
  assign _T_7159 = _T_2556 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26672.4]
  assign _T_7160 = _T_2816 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26673.4]
  assign _T_7162 = _T_7160 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26675.4]
  assign _T_7164 = _T_7154 + _T_7159; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26677.4]
  assign _T_7165 = _T_7164 - _T_7162; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26678.4]
  assign _T_7166 = $unsigned(_T_7165); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26679.4]
  assign _T_7167 = _T_7166[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26680.4]
  assign _T_7168 = _T_7162 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26682.4]
  assign _T_7170 = _T_7168 | _T_7154; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26684.4]
  assign _T_7172 = _T_7170 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26686.4]
  assign _T_7173 = _T_7172 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26687.4]
  assign _T_7174 = _T_7159 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26692.4]
  assign _T_7175 = _T_7154 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26693.4]
  assign _T_7176 = _T_7174 | _T_7175; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26694.4]
  assign _T_7178 = _T_7176 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26696.4]
  assign _T_7179 = _T_7178 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26697.4]
  assign _T_7190 = _T_2557 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26714.4]
  assign _T_7191 = _T_2817 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26715.4]
  assign _T_7193 = _T_7191 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26717.4]
  assign _T_7195 = _T_7185 + _T_7190; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26719.4]
  assign _T_7196 = _T_7195 - _T_7193; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26720.4]
  assign _T_7197 = $unsigned(_T_7196); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26721.4]
  assign _T_7198 = _T_7197[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26722.4]
  assign _T_7199 = _T_7193 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26724.4]
  assign _T_7201 = _T_7199 | _T_7185; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26726.4]
  assign _T_7203 = _T_7201 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26728.4]
  assign _T_7204 = _T_7203 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26729.4]
  assign _T_7205 = _T_7190 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26734.4]
  assign _T_7206 = _T_7185 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26735.4]
  assign _T_7207 = _T_7205 | _T_7206; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26736.4]
  assign _T_7209 = _T_7207 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26738.4]
  assign _T_7210 = _T_7209 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26739.4]
  assign _T_7221 = _T_2558 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26756.4]
  assign _T_7222 = _T_2818 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26757.4]
  assign _T_7224 = _T_7222 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26759.4]
  assign _T_7226 = _T_7216 + _T_7221; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26761.4]
  assign _T_7227 = _T_7226 - _T_7224; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26762.4]
  assign _T_7228 = $unsigned(_T_7227); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26763.4]
  assign _T_7229 = _T_7228[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26764.4]
  assign _T_7230 = _T_7224 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26766.4]
  assign _T_7232 = _T_7230 | _T_7216; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26768.4]
  assign _T_7234 = _T_7232 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26770.4]
  assign _T_7235 = _T_7234 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26771.4]
  assign _T_7236 = _T_7221 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26776.4]
  assign _T_7237 = _T_7216 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26777.4]
  assign _T_7238 = _T_7236 | _T_7237; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26778.4]
  assign _T_7240 = _T_7238 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26780.4]
  assign _T_7241 = _T_7240 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26781.4]
  assign _T_7252 = _T_2559 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26798.4]
  assign _T_7253 = _T_2819 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26799.4]
  assign _T_7255 = _T_7253 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26801.4]
  assign _T_7257 = _T_7247 + _T_7252; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26803.4]
  assign _T_7258 = _T_7257 - _T_7255; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26804.4]
  assign _T_7259 = $unsigned(_T_7258); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26805.4]
  assign _T_7260 = _T_7259[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26806.4]
  assign _T_7261 = _T_7255 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26808.4]
  assign _T_7263 = _T_7261 | _T_7247; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26810.4]
  assign _T_7265 = _T_7263 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26812.4]
  assign _T_7266 = _T_7265 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26813.4]
  assign _T_7267 = _T_7252 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26818.4]
  assign _T_7268 = _T_7247 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26819.4]
  assign _T_7269 = _T_7267 | _T_7268; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26820.4]
  assign _T_7271 = _T_7269 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26822.4]
  assign _T_7272 = _T_7271 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26823.4]
  assign _T_7283 = _T_2560 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26840.4]
  assign _T_7284 = _T_2820 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26841.4]
  assign _T_7286 = _T_7284 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26843.4]
  assign _T_7288 = _T_7278 + _T_7283; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26845.4]
  assign _T_7289 = _T_7288 - _T_7286; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26846.4]
  assign _T_7290 = $unsigned(_T_7289); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26847.4]
  assign _T_7291 = _T_7290[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26848.4]
  assign _T_7292 = _T_7286 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26850.4]
  assign _T_7294 = _T_7292 | _T_7278; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26852.4]
  assign _T_7296 = _T_7294 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26854.4]
  assign _T_7297 = _T_7296 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26855.4]
  assign _T_7298 = _T_7283 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26860.4]
  assign _T_7299 = _T_7278 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26861.4]
  assign _T_7300 = _T_7298 | _T_7299; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26862.4]
  assign _T_7302 = _T_7300 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26864.4]
  assign _T_7303 = _T_7302 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26865.4]
  assign _T_7314 = _T_2561 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26882.4]
  assign _T_7315 = _T_2821 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26883.4]
  assign _T_7317 = _T_7315 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26885.4]
  assign _T_7319 = _T_7309 + _T_7314; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26887.4]
  assign _T_7320 = _T_7319 - _T_7317; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26888.4]
  assign _T_7321 = $unsigned(_T_7320); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26889.4]
  assign _T_7322 = _T_7321[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26890.4]
  assign _T_7323 = _T_7317 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26892.4]
  assign _T_7325 = _T_7323 | _T_7309; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26894.4]
  assign _T_7327 = _T_7325 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26896.4]
  assign _T_7328 = _T_7327 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26897.4]
  assign _T_7329 = _T_7314 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26902.4]
  assign _T_7330 = _T_7309 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26903.4]
  assign _T_7331 = _T_7329 | _T_7330; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26904.4]
  assign _T_7333 = _T_7331 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26906.4]
  assign _T_7334 = _T_7333 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26907.4]
  assign _T_7345 = _T_2562 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26924.4]
  assign _T_7346 = _T_2822 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26925.4]
  assign _T_7348 = _T_7346 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26927.4]
  assign _T_7350 = _T_7340 + _T_7345; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26929.4]
  assign _T_7351 = _T_7350 - _T_7348; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26930.4]
  assign _T_7352 = $unsigned(_T_7351); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26931.4]
  assign _T_7353 = _T_7352[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26932.4]
  assign _T_7354 = _T_7348 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26934.4]
  assign _T_7356 = _T_7354 | _T_7340; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26936.4]
  assign _T_7358 = _T_7356 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26938.4]
  assign _T_7359 = _T_7358 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26939.4]
  assign _T_7360 = _T_7345 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26944.4]
  assign _T_7361 = _T_7340 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26945.4]
  assign _T_7362 = _T_7360 | _T_7361; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26946.4]
  assign _T_7364 = _T_7362 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26948.4]
  assign _T_7365 = _T_7364 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26949.4]
  assign _T_7376 = _T_2563 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@26966.4]
  assign _T_7377 = _T_2823 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@26967.4]
  assign _T_7379 = _T_7377 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@26969.4]
  assign _T_7381 = _T_7371 + _T_7376; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@26971.4]
  assign _T_7382 = _T_7381 - _T_7379; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26972.4]
  assign _T_7383 = $unsigned(_T_7382); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26973.4]
  assign _T_7384 = _T_7383[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@26974.4]
  assign _T_7385 = _T_7379 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@26976.4]
  assign _T_7387 = _T_7385 | _T_7371; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@26978.4]
  assign _T_7389 = _T_7387 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26980.4]
  assign _T_7390 = _T_7389 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26981.4]
  assign _T_7391 = _T_7376 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@26986.4]
  assign _T_7392 = _T_7371 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@26987.4]
  assign _T_7393 = _T_7391 | _T_7392; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@26988.4]
  assign _T_7395 = _T_7393 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26990.4]
  assign _T_7396 = _T_7395 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26991.4]
  assign _T_7407 = _T_2564 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27008.4]
  assign _T_7408 = _T_2824 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27009.4]
  assign _T_7410 = _T_7408 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27011.4]
  assign _T_7412 = _T_7402 + _T_7407; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27013.4]
  assign _T_7413 = _T_7412 - _T_7410; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27014.4]
  assign _T_7414 = $unsigned(_T_7413); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27015.4]
  assign _T_7415 = _T_7414[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27016.4]
  assign _T_7416 = _T_7410 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27018.4]
  assign _T_7418 = _T_7416 | _T_7402; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27020.4]
  assign _T_7420 = _T_7418 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27022.4]
  assign _T_7421 = _T_7420 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27023.4]
  assign _T_7422 = _T_7407 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27028.4]
  assign _T_7423 = _T_7402 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27029.4]
  assign _T_7424 = _T_7422 | _T_7423; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27030.4]
  assign _T_7426 = _T_7424 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27032.4]
  assign _T_7427 = _T_7426 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27033.4]
  assign _T_7438 = _T_2565 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27050.4]
  assign _T_7439 = _T_2825 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27051.4]
  assign _T_7441 = _T_7439 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27053.4]
  assign _T_7443 = _T_7433 + _T_7438; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27055.4]
  assign _T_7444 = _T_7443 - _T_7441; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27056.4]
  assign _T_7445 = $unsigned(_T_7444); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27057.4]
  assign _T_7446 = _T_7445[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27058.4]
  assign _T_7447 = _T_7441 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27060.4]
  assign _T_7449 = _T_7447 | _T_7433; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27062.4]
  assign _T_7451 = _T_7449 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27064.4]
  assign _T_7452 = _T_7451 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27065.4]
  assign _T_7453 = _T_7438 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27070.4]
  assign _T_7454 = _T_7433 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27071.4]
  assign _T_7455 = _T_7453 | _T_7454; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27072.4]
  assign _T_7457 = _T_7455 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27074.4]
  assign _T_7458 = _T_7457 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27075.4]
  assign _T_7469 = _T_2566 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27092.4]
  assign _T_7470 = _T_2826 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27093.4]
  assign _T_7472 = _T_7470 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27095.4]
  assign _T_7474 = _T_7464 + _T_7469; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27097.4]
  assign _T_7475 = _T_7474 - _T_7472; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27098.4]
  assign _T_7476 = $unsigned(_T_7475); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27099.4]
  assign _T_7477 = _T_7476[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27100.4]
  assign _T_7478 = _T_7472 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27102.4]
  assign _T_7480 = _T_7478 | _T_7464; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27104.4]
  assign _T_7482 = _T_7480 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27106.4]
  assign _T_7483 = _T_7482 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27107.4]
  assign _T_7484 = _T_7469 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27112.4]
  assign _T_7485 = _T_7464 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27113.4]
  assign _T_7486 = _T_7484 | _T_7485; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27114.4]
  assign _T_7488 = _T_7486 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27116.4]
  assign _T_7489 = _T_7488 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27117.4]
  assign _T_7500 = _T_2567 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27134.4]
  assign _T_7501 = _T_2827 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27135.4]
  assign _T_7503 = _T_7501 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27137.4]
  assign _T_7505 = _T_7495 + _T_7500; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27139.4]
  assign _T_7506 = _T_7505 - _T_7503; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27140.4]
  assign _T_7507 = $unsigned(_T_7506); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27141.4]
  assign _T_7508 = _T_7507[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27142.4]
  assign _T_7509 = _T_7503 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27144.4]
  assign _T_7511 = _T_7509 | _T_7495; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27146.4]
  assign _T_7513 = _T_7511 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27148.4]
  assign _T_7514 = _T_7513 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27149.4]
  assign _T_7515 = _T_7500 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27154.4]
  assign _T_7516 = _T_7495 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27155.4]
  assign _T_7517 = _T_7515 | _T_7516; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27156.4]
  assign _T_7519 = _T_7517 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27158.4]
  assign _T_7520 = _T_7519 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27159.4]
  assign _T_7531 = _T_2568 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27176.4]
  assign _T_7532 = _T_2828 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27177.4]
  assign _T_7534 = _T_7532 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27179.4]
  assign _T_7536 = _T_7526 + _T_7531; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27181.4]
  assign _T_7537 = _T_7536 - _T_7534; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27182.4]
  assign _T_7538 = $unsigned(_T_7537); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27183.4]
  assign _T_7539 = _T_7538[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27184.4]
  assign _T_7540 = _T_7534 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27186.4]
  assign _T_7542 = _T_7540 | _T_7526; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27188.4]
  assign _T_7544 = _T_7542 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27190.4]
  assign _T_7545 = _T_7544 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27191.4]
  assign _T_7546 = _T_7531 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27196.4]
  assign _T_7547 = _T_7526 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27197.4]
  assign _T_7548 = _T_7546 | _T_7547; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27198.4]
  assign _T_7550 = _T_7548 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27200.4]
  assign _T_7551 = _T_7550 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27201.4]
  assign _T_7562 = _T_2569 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27218.4]
  assign _T_7563 = _T_2829 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27219.4]
  assign _T_7565 = _T_7563 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27221.4]
  assign _T_7567 = _T_7557 + _T_7562; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27223.4]
  assign _T_7568 = _T_7567 - _T_7565; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27224.4]
  assign _T_7569 = $unsigned(_T_7568); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27225.4]
  assign _T_7570 = _T_7569[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27226.4]
  assign _T_7571 = _T_7565 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27228.4]
  assign _T_7573 = _T_7571 | _T_7557; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27230.4]
  assign _T_7575 = _T_7573 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27232.4]
  assign _T_7576 = _T_7575 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27233.4]
  assign _T_7577 = _T_7562 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27238.4]
  assign _T_7578 = _T_7557 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27239.4]
  assign _T_7579 = _T_7577 | _T_7578; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27240.4]
  assign _T_7581 = _T_7579 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27242.4]
  assign _T_7582 = _T_7581 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27243.4]
  assign _T_7593 = _T_2570 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27260.4]
  assign _T_7594 = _T_2830 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27261.4]
  assign _T_7596 = _T_7594 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27263.4]
  assign _T_7598 = _T_7588 + _T_7593; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27265.4]
  assign _T_7599 = _T_7598 - _T_7596; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27266.4]
  assign _T_7600 = $unsigned(_T_7599); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27267.4]
  assign _T_7601 = _T_7600[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27268.4]
  assign _T_7602 = _T_7596 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27270.4]
  assign _T_7604 = _T_7602 | _T_7588; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27272.4]
  assign _T_7606 = _T_7604 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27274.4]
  assign _T_7607 = _T_7606 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27275.4]
  assign _T_7608 = _T_7593 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27280.4]
  assign _T_7609 = _T_7588 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27281.4]
  assign _T_7610 = _T_7608 | _T_7609; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27282.4]
  assign _T_7612 = _T_7610 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27284.4]
  assign _T_7613 = _T_7612 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27285.4]
  assign _T_7624 = _T_2571 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27302.4]
  assign _T_7625 = _T_2831 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27303.4]
  assign _T_7627 = _T_7625 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27305.4]
  assign _T_7629 = _T_7619 + _T_7624; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27307.4]
  assign _T_7630 = _T_7629 - _T_7627; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27308.4]
  assign _T_7631 = $unsigned(_T_7630); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27309.4]
  assign _T_7632 = _T_7631[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27310.4]
  assign _T_7633 = _T_7627 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27312.4]
  assign _T_7635 = _T_7633 | _T_7619; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27314.4]
  assign _T_7637 = _T_7635 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27316.4]
  assign _T_7638 = _T_7637 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27317.4]
  assign _T_7639 = _T_7624 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27322.4]
  assign _T_7640 = _T_7619 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27323.4]
  assign _T_7641 = _T_7639 | _T_7640; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27324.4]
  assign _T_7643 = _T_7641 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27326.4]
  assign _T_7644 = _T_7643 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27327.4]
  assign _T_7655 = _T_2572 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27344.4]
  assign _T_7656 = _T_2832 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27345.4]
  assign _T_7658 = _T_7656 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27347.4]
  assign _T_7660 = _T_7650 + _T_7655; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27349.4]
  assign _T_7661 = _T_7660 - _T_7658; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27350.4]
  assign _T_7662 = $unsigned(_T_7661); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27351.4]
  assign _T_7663 = _T_7662[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27352.4]
  assign _T_7664 = _T_7658 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27354.4]
  assign _T_7666 = _T_7664 | _T_7650; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27356.4]
  assign _T_7668 = _T_7666 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27358.4]
  assign _T_7669 = _T_7668 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27359.4]
  assign _T_7670 = _T_7655 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27364.4]
  assign _T_7671 = _T_7650 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27365.4]
  assign _T_7672 = _T_7670 | _T_7671; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27366.4]
  assign _T_7674 = _T_7672 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27368.4]
  assign _T_7675 = _T_7674 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27369.4]
  assign _T_7686 = _T_2573 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27386.4]
  assign _T_7687 = _T_2833 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27387.4]
  assign _T_7689 = _T_7687 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27389.4]
  assign _T_7691 = _T_7681 + _T_7686; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27391.4]
  assign _T_7692 = _T_7691 - _T_7689; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27392.4]
  assign _T_7693 = $unsigned(_T_7692); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27393.4]
  assign _T_7694 = _T_7693[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27394.4]
  assign _T_7695 = _T_7689 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27396.4]
  assign _T_7697 = _T_7695 | _T_7681; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27398.4]
  assign _T_7699 = _T_7697 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27400.4]
  assign _T_7700 = _T_7699 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27401.4]
  assign _T_7701 = _T_7686 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27406.4]
  assign _T_7702 = _T_7681 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27407.4]
  assign _T_7703 = _T_7701 | _T_7702; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27408.4]
  assign _T_7705 = _T_7703 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27410.4]
  assign _T_7706 = _T_7705 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27411.4]
  assign _T_7717 = _T_2574 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27428.4]
  assign _T_7718 = _T_2834 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27429.4]
  assign _T_7720 = _T_7718 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27431.4]
  assign _T_7722 = _T_7712 + _T_7717; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27433.4]
  assign _T_7723 = _T_7722 - _T_7720; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27434.4]
  assign _T_7724 = $unsigned(_T_7723); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27435.4]
  assign _T_7725 = _T_7724[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27436.4]
  assign _T_7726 = _T_7720 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27438.4]
  assign _T_7728 = _T_7726 | _T_7712; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27440.4]
  assign _T_7730 = _T_7728 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27442.4]
  assign _T_7731 = _T_7730 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27443.4]
  assign _T_7732 = _T_7717 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27448.4]
  assign _T_7733 = _T_7712 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27449.4]
  assign _T_7734 = _T_7732 | _T_7733; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27450.4]
  assign _T_7736 = _T_7734 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27452.4]
  assign _T_7737 = _T_7736 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27453.4]
  assign _T_7748 = _T_2575 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27470.4]
  assign _T_7749 = _T_2835 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27471.4]
  assign _T_7751 = _T_7749 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27473.4]
  assign _T_7753 = _T_7743 + _T_7748; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27475.4]
  assign _T_7754 = _T_7753 - _T_7751; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27476.4]
  assign _T_7755 = $unsigned(_T_7754); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27477.4]
  assign _T_7756 = _T_7755[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27478.4]
  assign _T_7757 = _T_7751 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27480.4]
  assign _T_7759 = _T_7757 | _T_7743; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27482.4]
  assign _T_7761 = _T_7759 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27484.4]
  assign _T_7762 = _T_7761 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27485.4]
  assign _T_7763 = _T_7748 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27490.4]
  assign _T_7764 = _T_7743 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27491.4]
  assign _T_7765 = _T_7763 | _T_7764; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27492.4]
  assign _T_7767 = _T_7765 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27494.4]
  assign _T_7768 = _T_7767 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27495.4]
  assign _T_7779 = _T_2576 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27512.4]
  assign _T_7780 = _T_2836 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27513.4]
  assign _T_7782 = _T_7780 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27515.4]
  assign _T_7784 = _T_7774 + _T_7779; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27517.4]
  assign _T_7785 = _T_7784 - _T_7782; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27518.4]
  assign _T_7786 = $unsigned(_T_7785); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27519.4]
  assign _T_7787 = _T_7786[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27520.4]
  assign _T_7788 = _T_7782 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27522.4]
  assign _T_7790 = _T_7788 | _T_7774; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27524.4]
  assign _T_7792 = _T_7790 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27526.4]
  assign _T_7793 = _T_7792 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27527.4]
  assign _T_7794 = _T_7779 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27532.4]
  assign _T_7795 = _T_7774 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27533.4]
  assign _T_7796 = _T_7794 | _T_7795; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27534.4]
  assign _T_7798 = _T_7796 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27536.4]
  assign _T_7799 = _T_7798 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27537.4]
  assign _T_7810 = _T_2577 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27554.4]
  assign _T_7811 = _T_2837 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27555.4]
  assign _T_7813 = _T_7811 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27557.4]
  assign _T_7815 = _T_7805 + _T_7810; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27559.4]
  assign _T_7816 = _T_7815 - _T_7813; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27560.4]
  assign _T_7817 = $unsigned(_T_7816); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27561.4]
  assign _T_7818 = _T_7817[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27562.4]
  assign _T_7819 = _T_7813 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27564.4]
  assign _T_7821 = _T_7819 | _T_7805; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27566.4]
  assign _T_7823 = _T_7821 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27568.4]
  assign _T_7824 = _T_7823 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27569.4]
  assign _T_7825 = _T_7810 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27574.4]
  assign _T_7826 = _T_7805 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27575.4]
  assign _T_7827 = _T_7825 | _T_7826; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27576.4]
  assign _T_7829 = _T_7827 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27578.4]
  assign _T_7830 = _T_7829 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27579.4]
  assign _T_7841 = _T_2578 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27596.4]
  assign _T_7842 = _T_2838 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27597.4]
  assign _T_7844 = _T_7842 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27599.4]
  assign _T_7846 = _T_7836 + _T_7841; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27601.4]
  assign _T_7847 = _T_7846 - _T_7844; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27602.4]
  assign _T_7848 = $unsigned(_T_7847); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27603.4]
  assign _T_7849 = _T_7848[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27604.4]
  assign _T_7850 = _T_7844 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27606.4]
  assign _T_7852 = _T_7850 | _T_7836; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27608.4]
  assign _T_7854 = _T_7852 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27610.4]
  assign _T_7855 = _T_7854 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27611.4]
  assign _T_7856 = _T_7841 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27616.4]
  assign _T_7857 = _T_7836 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27617.4]
  assign _T_7858 = _T_7856 | _T_7857; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27618.4]
  assign _T_7860 = _T_7858 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27620.4]
  assign _T_7861 = _T_7860 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27621.4]
  assign _T_7872 = _T_2579 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27638.4]
  assign _T_7873 = _T_2839 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27639.4]
  assign _T_7875 = _T_7873 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27641.4]
  assign _T_7877 = _T_7867 + _T_7872; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27643.4]
  assign _T_7878 = _T_7877 - _T_7875; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27644.4]
  assign _T_7879 = $unsigned(_T_7878); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27645.4]
  assign _T_7880 = _T_7879[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27646.4]
  assign _T_7881 = _T_7875 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27648.4]
  assign _T_7883 = _T_7881 | _T_7867; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27650.4]
  assign _T_7885 = _T_7883 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27652.4]
  assign _T_7886 = _T_7885 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27653.4]
  assign _T_7887 = _T_7872 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27658.4]
  assign _T_7888 = _T_7867 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27659.4]
  assign _T_7889 = _T_7887 | _T_7888; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27660.4]
  assign _T_7891 = _T_7889 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27662.4]
  assign _T_7892 = _T_7891 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27663.4]
  assign _T_7903 = _T_2580 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27680.4]
  assign _T_7904 = _T_2840 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27681.4]
  assign _T_7906 = _T_7904 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27683.4]
  assign _T_7908 = _T_7898 + _T_7903; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27685.4]
  assign _T_7909 = _T_7908 - _T_7906; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27686.4]
  assign _T_7910 = $unsigned(_T_7909); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27687.4]
  assign _T_7911 = _T_7910[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27688.4]
  assign _T_7912 = _T_7906 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27690.4]
  assign _T_7914 = _T_7912 | _T_7898; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27692.4]
  assign _T_7916 = _T_7914 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27694.4]
  assign _T_7917 = _T_7916 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27695.4]
  assign _T_7918 = _T_7903 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27700.4]
  assign _T_7919 = _T_7898 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27701.4]
  assign _T_7920 = _T_7918 | _T_7919; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27702.4]
  assign _T_7922 = _T_7920 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27704.4]
  assign _T_7923 = _T_7922 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27705.4]
  assign _T_7934 = _T_2581 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27722.4]
  assign _T_7935 = _T_2841 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27723.4]
  assign _T_7937 = _T_7935 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27725.4]
  assign _T_7939 = _T_7929 + _T_7934; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27727.4]
  assign _T_7940 = _T_7939 - _T_7937; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27728.4]
  assign _T_7941 = $unsigned(_T_7940); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27729.4]
  assign _T_7942 = _T_7941[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27730.4]
  assign _T_7943 = _T_7937 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27732.4]
  assign _T_7945 = _T_7943 | _T_7929; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27734.4]
  assign _T_7947 = _T_7945 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27736.4]
  assign _T_7948 = _T_7947 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27737.4]
  assign _T_7949 = _T_7934 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27742.4]
  assign _T_7950 = _T_7929 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27743.4]
  assign _T_7951 = _T_7949 | _T_7950; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27744.4]
  assign _T_7953 = _T_7951 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27746.4]
  assign _T_7954 = _T_7953 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27747.4]
  assign _T_7965 = _T_2582 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27764.4]
  assign _T_7966 = _T_2842 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27765.4]
  assign _T_7968 = _T_7966 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27767.4]
  assign _T_7970 = _T_7960 + _T_7965; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27769.4]
  assign _T_7971 = _T_7970 - _T_7968; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27770.4]
  assign _T_7972 = $unsigned(_T_7971); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27771.4]
  assign _T_7973 = _T_7972[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27772.4]
  assign _T_7974 = _T_7968 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27774.4]
  assign _T_7976 = _T_7974 | _T_7960; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27776.4]
  assign _T_7978 = _T_7976 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27778.4]
  assign _T_7979 = _T_7978 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27779.4]
  assign _T_7980 = _T_7965 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27784.4]
  assign _T_7981 = _T_7960 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27785.4]
  assign _T_7982 = _T_7980 | _T_7981; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27786.4]
  assign _T_7984 = _T_7982 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27788.4]
  assign _T_7985 = _T_7984 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27789.4]
  assign _T_7996 = _T_2583 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27806.4]
  assign _T_7997 = _T_2843 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27807.4]
  assign _T_7999 = _T_7997 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27809.4]
  assign _T_8001 = _T_7991 + _T_7996; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27811.4]
  assign _T_8002 = _T_8001 - _T_7999; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27812.4]
  assign _T_8003 = $unsigned(_T_8002); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27813.4]
  assign _T_8004 = _T_8003[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27814.4]
  assign _T_8005 = _T_7999 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27816.4]
  assign _T_8007 = _T_8005 | _T_7991; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27818.4]
  assign _T_8009 = _T_8007 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27820.4]
  assign _T_8010 = _T_8009 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27821.4]
  assign _T_8011 = _T_7996 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27826.4]
  assign _T_8012 = _T_7991 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27827.4]
  assign _T_8013 = _T_8011 | _T_8012; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27828.4]
  assign _T_8015 = _T_8013 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27830.4]
  assign _T_8016 = _T_8015 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27831.4]
  assign _T_8027 = _T_2584 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27848.4]
  assign _T_8028 = _T_2844 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27849.4]
  assign _T_8030 = _T_8028 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27851.4]
  assign _T_8032 = _T_8022 + _T_8027; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27853.4]
  assign _T_8033 = _T_8032 - _T_8030; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27854.4]
  assign _T_8034 = $unsigned(_T_8033); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27855.4]
  assign _T_8035 = _T_8034[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27856.4]
  assign _T_8036 = _T_8030 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27858.4]
  assign _T_8038 = _T_8036 | _T_8022; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27860.4]
  assign _T_8040 = _T_8038 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27862.4]
  assign _T_8041 = _T_8040 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27863.4]
  assign _T_8042 = _T_8027 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27868.4]
  assign _T_8043 = _T_8022 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27869.4]
  assign _T_8044 = _T_8042 | _T_8043; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27870.4]
  assign _T_8046 = _T_8044 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27872.4]
  assign _T_8047 = _T_8046 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27873.4]
  assign _T_8058 = _T_2585 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27890.4]
  assign _T_8059 = _T_2845 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27891.4]
  assign _T_8061 = _T_8059 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27893.4]
  assign _T_8063 = _T_8053 + _T_8058; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27895.4]
  assign _T_8064 = _T_8063 - _T_8061; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27896.4]
  assign _T_8065 = $unsigned(_T_8064); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27897.4]
  assign _T_8066 = _T_8065[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27898.4]
  assign _T_8067 = _T_8061 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27900.4]
  assign _T_8069 = _T_8067 | _T_8053; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27902.4]
  assign _T_8071 = _T_8069 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27904.4]
  assign _T_8072 = _T_8071 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27905.4]
  assign _T_8073 = _T_8058 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27910.4]
  assign _T_8074 = _T_8053 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27911.4]
  assign _T_8075 = _T_8073 | _T_8074; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27912.4]
  assign _T_8077 = _T_8075 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27914.4]
  assign _T_8078 = _T_8077 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27915.4]
  assign _T_8089 = _T_2586 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27932.4]
  assign _T_8090 = _T_2846 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27933.4]
  assign _T_8092 = _T_8090 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27935.4]
  assign _T_8094 = _T_8084 + _T_8089; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27937.4]
  assign _T_8095 = _T_8094 - _T_8092; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27938.4]
  assign _T_8096 = $unsigned(_T_8095); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27939.4]
  assign _T_8097 = _T_8096[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27940.4]
  assign _T_8098 = _T_8092 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27942.4]
  assign _T_8100 = _T_8098 | _T_8084; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27944.4]
  assign _T_8102 = _T_8100 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27946.4]
  assign _T_8103 = _T_8102 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27947.4]
  assign _T_8104 = _T_8089 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27952.4]
  assign _T_8105 = _T_8084 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27953.4]
  assign _T_8106 = _T_8104 | _T_8105; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27954.4]
  assign _T_8108 = _T_8106 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27956.4]
  assign _T_8109 = _T_8108 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27957.4]
  assign _T_8120 = _T_2587 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@27974.4]
  assign _T_8121 = _T_2847 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@27975.4]
  assign _T_8123 = _T_8121 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@27977.4]
  assign _T_8125 = _T_8115 + _T_8120; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@27979.4]
  assign _T_8126 = _T_8125 - _T_8123; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27980.4]
  assign _T_8127 = $unsigned(_T_8126); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27981.4]
  assign _T_8128 = _T_8127[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@27982.4]
  assign _T_8129 = _T_8123 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@27984.4]
  assign _T_8131 = _T_8129 | _T_8115; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@27986.4]
  assign _T_8133 = _T_8131 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27988.4]
  assign _T_8134 = _T_8133 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27989.4]
  assign _T_8135 = _T_8120 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@27994.4]
  assign _T_8136 = _T_8115 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@27995.4]
  assign _T_8137 = _T_8135 | _T_8136; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@27996.4]
  assign _T_8139 = _T_8137 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27998.4]
  assign _T_8140 = _T_8139 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27999.4]
  assign _T_8151 = _T_2588 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28016.4]
  assign _T_8152 = _T_2848 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28017.4]
  assign _T_8154 = _T_8152 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28019.4]
  assign _T_8156 = _T_8146 + _T_8151; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28021.4]
  assign _T_8157 = _T_8156 - _T_8154; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28022.4]
  assign _T_8158 = $unsigned(_T_8157); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28023.4]
  assign _T_8159 = _T_8158[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28024.4]
  assign _T_8160 = _T_8154 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28026.4]
  assign _T_8162 = _T_8160 | _T_8146; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28028.4]
  assign _T_8164 = _T_8162 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28030.4]
  assign _T_8165 = _T_8164 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28031.4]
  assign _T_8166 = _T_8151 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28036.4]
  assign _T_8167 = _T_8146 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28037.4]
  assign _T_8168 = _T_8166 | _T_8167; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28038.4]
  assign _T_8170 = _T_8168 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28040.4]
  assign _T_8171 = _T_8170 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28041.4]
  assign _T_8182 = _T_2589 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28058.4]
  assign _T_8183 = _T_2849 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28059.4]
  assign _T_8185 = _T_8183 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28061.4]
  assign _T_8187 = _T_8177 + _T_8182; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28063.4]
  assign _T_8188 = _T_8187 - _T_8185; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28064.4]
  assign _T_8189 = $unsigned(_T_8188); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28065.4]
  assign _T_8190 = _T_8189[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28066.4]
  assign _T_8191 = _T_8185 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28068.4]
  assign _T_8193 = _T_8191 | _T_8177; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28070.4]
  assign _T_8195 = _T_8193 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28072.4]
  assign _T_8196 = _T_8195 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28073.4]
  assign _T_8197 = _T_8182 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28078.4]
  assign _T_8198 = _T_8177 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28079.4]
  assign _T_8199 = _T_8197 | _T_8198; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28080.4]
  assign _T_8201 = _T_8199 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28082.4]
  assign _T_8202 = _T_8201 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28083.4]
  assign _T_8213 = _T_2590 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28100.4]
  assign _T_8214 = _T_2850 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28101.4]
  assign _T_8216 = _T_8214 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28103.4]
  assign _T_8218 = _T_8208 + _T_8213; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28105.4]
  assign _T_8219 = _T_8218 - _T_8216; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28106.4]
  assign _T_8220 = $unsigned(_T_8219); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28107.4]
  assign _T_8221 = _T_8220[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28108.4]
  assign _T_8222 = _T_8216 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28110.4]
  assign _T_8224 = _T_8222 | _T_8208; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28112.4]
  assign _T_8226 = _T_8224 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28114.4]
  assign _T_8227 = _T_8226 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28115.4]
  assign _T_8228 = _T_8213 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28120.4]
  assign _T_8229 = _T_8208 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28121.4]
  assign _T_8230 = _T_8228 | _T_8229; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28122.4]
  assign _T_8232 = _T_8230 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28124.4]
  assign _T_8233 = _T_8232 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28125.4]
  assign _T_8244 = _T_2591 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28142.4]
  assign _T_8245 = _T_2851 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28143.4]
  assign _T_8247 = _T_8245 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28145.4]
  assign _T_8249 = _T_8239 + _T_8244; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28147.4]
  assign _T_8250 = _T_8249 - _T_8247; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28148.4]
  assign _T_8251 = $unsigned(_T_8250); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28149.4]
  assign _T_8252 = _T_8251[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28150.4]
  assign _T_8253 = _T_8247 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28152.4]
  assign _T_8255 = _T_8253 | _T_8239; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28154.4]
  assign _T_8257 = _T_8255 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28156.4]
  assign _T_8258 = _T_8257 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28157.4]
  assign _T_8259 = _T_8244 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28162.4]
  assign _T_8260 = _T_8239 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28163.4]
  assign _T_8261 = _T_8259 | _T_8260; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28164.4]
  assign _T_8263 = _T_8261 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28166.4]
  assign _T_8264 = _T_8263 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28167.4]
  assign _T_8275 = _T_2592 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28184.4]
  assign _T_8276 = _T_2852 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28185.4]
  assign _T_8278 = _T_8276 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28187.4]
  assign _T_8280 = _T_8270 + _T_8275; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28189.4]
  assign _T_8281 = _T_8280 - _T_8278; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28190.4]
  assign _T_8282 = $unsigned(_T_8281); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28191.4]
  assign _T_8283 = _T_8282[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28192.4]
  assign _T_8284 = _T_8278 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28194.4]
  assign _T_8286 = _T_8284 | _T_8270; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28196.4]
  assign _T_8288 = _T_8286 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28198.4]
  assign _T_8289 = _T_8288 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28199.4]
  assign _T_8290 = _T_8275 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28204.4]
  assign _T_8291 = _T_8270 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28205.4]
  assign _T_8292 = _T_8290 | _T_8291; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28206.4]
  assign _T_8294 = _T_8292 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28208.4]
  assign _T_8295 = _T_8294 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28209.4]
  assign _T_8306 = _T_2593 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28226.4]
  assign _T_8307 = _T_2853 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28227.4]
  assign _T_8309 = _T_8307 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28229.4]
  assign _T_8311 = _T_8301 + _T_8306; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28231.4]
  assign _T_8312 = _T_8311 - _T_8309; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28232.4]
  assign _T_8313 = $unsigned(_T_8312); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28233.4]
  assign _T_8314 = _T_8313[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28234.4]
  assign _T_8315 = _T_8309 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28236.4]
  assign _T_8317 = _T_8315 | _T_8301; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28238.4]
  assign _T_8319 = _T_8317 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28240.4]
  assign _T_8320 = _T_8319 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28241.4]
  assign _T_8321 = _T_8306 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28246.4]
  assign _T_8322 = _T_8301 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28247.4]
  assign _T_8323 = _T_8321 | _T_8322; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28248.4]
  assign _T_8325 = _T_8323 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28250.4]
  assign _T_8326 = _T_8325 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28251.4]
  assign _T_8337 = _T_2594 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28268.4]
  assign _T_8338 = _T_2854 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28269.4]
  assign _T_8340 = _T_8338 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28271.4]
  assign _T_8342 = _T_8332 + _T_8337; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28273.4]
  assign _T_8343 = _T_8342 - _T_8340; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28274.4]
  assign _T_8344 = $unsigned(_T_8343); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28275.4]
  assign _T_8345 = _T_8344[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28276.4]
  assign _T_8346 = _T_8340 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28278.4]
  assign _T_8348 = _T_8346 | _T_8332; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28280.4]
  assign _T_8350 = _T_8348 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28282.4]
  assign _T_8351 = _T_8350 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28283.4]
  assign _T_8352 = _T_8337 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28288.4]
  assign _T_8353 = _T_8332 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28289.4]
  assign _T_8354 = _T_8352 | _T_8353; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28290.4]
  assign _T_8356 = _T_8354 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28292.4]
  assign _T_8357 = _T_8356 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28293.4]
  assign _T_8368 = _T_2595 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28310.4]
  assign _T_8369 = _T_2855 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28311.4]
  assign _T_8371 = _T_8369 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28313.4]
  assign _T_8373 = _T_8363 + _T_8368; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28315.4]
  assign _T_8374 = _T_8373 - _T_8371; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28316.4]
  assign _T_8375 = $unsigned(_T_8374); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28317.4]
  assign _T_8376 = _T_8375[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28318.4]
  assign _T_8377 = _T_8371 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28320.4]
  assign _T_8379 = _T_8377 | _T_8363; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28322.4]
  assign _T_8381 = _T_8379 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28324.4]
  assign _T_8382 = _T_8381 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28325.4]
  assign _T_8383 = _T_8368 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28330.4]
  assign _T_8384 = _T_8363 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28331.4]
  assign _T_8385 = _T_8383 | _T_8384; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28332.4]
  assign _T_8387 = _T_8385 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28334.4]
  assign _T_8388 = _T_8387 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28335.4]
  assign _T_8399 = _T_2596 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28352.4]
  assign _T_8400 = _T_2856 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28353.4]
  assign _T_8402 = _T_8400 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28355.4]
  assign _T_8404 = _T_8394 + _T_8399; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28357.4]
  assign _T_8405 = _T_8404 - _T_8402; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28358.4]
  assign _T_8406 = $unsigned(_T_8405); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28359.4]
  assign _T_8407 = _T_8406[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28360.4]
  assign _T_8408 = _T_8402 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28362.4]
  assign _T_8410 = _T_8408 | _T_8394; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28364.4]
  assign _T_8412 = _T_8410 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28366.4]
  assign _T_8413 = _T_8412 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28367.4]
  assign _T_8414 = _T_8399 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28372.4]
  assign _T_8415 = _T_8394 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28373.4]
  assign _T_8416 = _T_8414 | _T_8415; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28374.4]
  assign _T_8418 = _T_8416 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28376.4]
  assign _T_8419 = _T_8418 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28377.4]
  assign _T_8430 = _T_2597 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28394.4]
  assign _T_8431 = _T_2857 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28395.4]
  assign _T_8433 = _T_8431 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28397.4]
  assign _T_8435 = _T_8425 + _T_8430; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28399.4]
  assign _T_8436 = _T_8435 - _T_8433; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28400.4]
  assign _T_8437 = $unsigned(_T_8436); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28401.4]
  assign _T_8438 = _T_8437[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28402.4]
  assign _T_8439 = _T_8433 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28404.4]
  assign _T_8441 = _T_8439 | _T_8425; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28406.4]
  assign _T_8443 = _T_8441 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28408.4]
  assign _T_8444 = _T_8443 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28409.4]
  assign _T_8445 = _T_8430 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28414.4]
  assign _T_8446 = _T_8425 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28415.4]
  assign _T_8447 = _T_8445 | _T_8446; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28416.4]
  assign _T_8449 = _T_8447 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28418.4]
  assign _T_8450 = _T_8449 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28419.4]
  assign _T_8461 = _T_2598 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28436.4]
  assign _T_8462 = _T_2858 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28437.4]
  assign _T_8464 = _T_8462 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28439.4]
  assign _T_8466 = _T_8456 + _T_8461; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28441.4]
  assign _T_8467 = _T_8466 - _T_8464; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28442.4]
  assign _T_8468 = $unsigned(_T_8467); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28443.4]
  assign _T_8469 = _T_8468[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28444.4]
  assign _T_8470 = _T_8464 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28446.4]
  assign _T_8472 = _T_8470 | _T_8456; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28448.4]
  assign _T_8474 = _T_8472 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28450.4]
  assign _T_8475 = _T_8474 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28451.4]
  assign _T_8476 = _T_8461 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28456.4]
  assign _T_8477 = _T_8456 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28457.4]
  assign _T_8478 = _T_8476 | _T_8477; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28458.4]
  assign _T_8480 = _T_8478 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28460.4]
  assign _T_8481 = _T_8480 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28461.4]
  assign _T_8492 = _T_2599 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28478.4]
  assign _T_8493 = _T_2859 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28479.4]
  assign _T_8495 = _T_8493 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28481.4]
  assign _T_8497 = _T_8487 + _T_8492; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28483.4]
  assign _T_8498 = _T_8497 - _T_8495; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28484.4]
  assign _T_8499 = $unsigned(_T_8498); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28485.4]
  assign _T_8500 = _T_8499[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28486.4]
  assign _T_8501 = _T_8495 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28488.4]
  assign _T_8503 = _T_8501 | _T_8487; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28490.4]
  assign _T_8505 = _T_8503 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28492.4]
  assign _T_8506 = _T_8505 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28493.4]
  assign _T_8507 = _T_8492 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28498.4]
  assign _T_8508 = _T_8487 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28499.4]
  assign _T_8509 = _T_8507 | _T_8508; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28500.4]
  assign _T_8511 = _T_8509 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28502.4]
  assign _T_8512 = _T_8511 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28503.4]
  assign _T_8523 = _T_2600 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28520.4]
  assign _T_8524 = _T_2860 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28521.4]
  assign _T_8526 = _T_8524 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28523.4]
  assign _T_8528 = _T_8518 + _T_8523; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28525.4]
  assign _T_8529 = _T_8528 - _T_8526; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28526.4]
  assign _T_8530 = $unsigned(_T_8529); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28527.4]
  assign _T_8531 = _T_8530[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28528.4]
  assign _T_8532 = _T_8526 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28530.4]
  assign _T_8534 = _T_8532 | _T_8518; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28532.4]
  assign _T_8536 = _T_8534 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28534.4]
  assign _T_8537 = _T_8536 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28535.4]
  assign _T_8538 = _T_8523 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28540.4]
  assign _T_8539 = _T_8518 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28541.4]
  assign _T_8540 = _T_8538 | _T_8539; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28542.4]
  assign _T_8542 = _T_8540 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28544.4]
  assign _T_8543 = _T_8542 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28545.4]
  assign _T_8554 = _T_2601 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28562.4]
  assign _T_8555 = _T_2861 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28563.4]
  assign _T_8557 = _T_8555 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28565.4]
  assign _T_8559 = _T_8549 + _T_8554; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28567.4]
  assign _T_8560 = _T_8559 - _T_8557; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28568.4]
  assign _T_8561 = $unsigned(_T_8560); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28569.4]
  assign _T_8562 = _T_8561[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28570.4]
  assign _T_8563 = _T_8557 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28572.4]
  assign _T_8565 = _T_8563 | _T_8549; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28574.4]
  assign _T_8567 = _T_8565 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28576.4]
  assign _T_8568 = _T_8567 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28577.4]
  assign _T_8569 = _T_8554 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28582.4]
  assign _T_8570 = _T_8549 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28583.4]
  assign _T_8571 = _T_8569 | _T_8570; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28584.4]
  assign _T_8573 = _T_8571 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28586.4]
  assign _T_8574 = _T_8573 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28587.4]
  assign _T_8585 = _T_2602 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28604.4]
  assign _T_8586 = _T_2862 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28605.4]
  assign _T_8588 = _T_8586 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28607.4]
  assign _T_8590 = _T_8580 + _T_8585; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28609.4]
  assign _T_8591 = _T_8590 - _T_8588; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28610.4]
  assign _T_8592 = $unsigned(_T_8591); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28611.4]
  assign _T_8593 = _T_8592[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28612.4]
  assign _T_8594 = _T_8588 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28614.4]
  assign _T_8596 = _T_8594 | _T_8580; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28616.4]
  assign _T_8598 = _T_8596 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28618.4]
  assign _T_8599 = _T_8598 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28619.4]
  assign _T_8600 = _T_8585 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28624.4]
  assign _T_8601 = _T_8580 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28625.4]
  assign _T_8602 = _T_8600 | _T_8601; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28626.4]
  assign _T_8604 = _T_8602 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28628.4]
  assign _T_8605 = _T_8604 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28629.4]
  assign _T_8616 = _T_2603 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28646.4]
  assign _T_8617 = _T_2863 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28647.4]
  assign _T_8619 = _T_8617 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28649.4]
  assign _T_8621 = _T_8611 + _T_8616; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28651.4]
  assign _T_8622 = _T_8621 - _T_8619; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28652.4]
  assign _T_8623 = $unsigned(_T_8622); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28653.4]
  assign _T_8624 = _T_8623[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28654.4]
  assign _T_8625 = _T_8619 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28656.4]
  assign _T_8627 = _T_8625 | _T_8611; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28658.4]
  assign _T_8629 = _T_8627 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28660.4]
  assign _T_8630 = _T_8629 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28661.4]
  assign _T_8631 = _T_8616 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28666.4]
  assign _T_8632 = _T_8611 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28667.4]
  assign _T_8633 = _T_8631 | _T_8632; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28668.4]
  assign _T_8635 = _T_8633 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28670.4]
  assign _T_8636 = _T_8635 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28671.4]
  assign _T_8647 = _T_2604 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28688.4]
  assign _T_8648 = _T_2864 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28689.4]
  assign _T_8650 = _T_8648 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28691.4]
  assign _T_8652 = _T_8642 + _T_8647; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28693.4]
  assign _T_8653 = _T_8652 - _T_8650; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28694.4]
  assign _T_8654 = $unsigned(_T_8653); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28695.4]
  assign _T_8655 = _T_8654[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28696.4]
  assign _T_8656 = _T_8650 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28698.4]
  assign _T_8658 = _T_8656 | _T_8642; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28700.4]
  assign _T_8660 = _T_8658 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28702.4]
  assign _T_8661 = _T_8660 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28703.4]
  assign _T_8662 = _T_8647 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28708.4]
  assign _T_8663 = _T_8642 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28709.4]
  assign _T_8664 = _T_8662 | _T_8663; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28710.4]
  assign _T_8666 = _T_8664 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28712.4]
  assign _T_8667 = _T_8666 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28713.4]
  assign _T_8678 = _T_2605 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28730.4]
  assign _T_8679 = _T_2865 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28731.4]
  assign _T_8681 = _T_8679 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28733.4]
  assign _T_8683 = _T_8673 + _T_8678; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28735.4]
  assign _T_8684 = _T_8683 - _T_8681; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28736.4]
  assign _T_8685 = $unsigned(_T_8684); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28737.4]
  assign _T_8686 = _T_8685[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28738.4]
  assign _T_8687 = _T_8681 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28740.4]
  assign _T_8689 = _T_8687 | _T_8673; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28742.4]
  assign _T_8691 = _T_8689 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28744.4]
  assign _T_8692 = _T_8691 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28745.4]
  assign _T_8693 = _T_8678 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28750.4]
  assign _T_8694 = _T_8673 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28751.4]
  assign _T_8695 = _T_8693 | _T_8694; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28752.4]
  assign _T_8697 = _T_8695 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28754.4]
  assign _T_8698 = _T_8697 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28755.4]
  assign _T_8709 = _T_2606 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28772.4]
  assign _T_8710 = _T_2866 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28773.4]
  assign _T_8712 = _T_8710 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28775.4]
  assign _T_8714 = _T_8704 + _T_8709; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28777.4]
  assign _T_8715 = _T_8714 - _T_8712; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28778.4]
  assign _T_8716 = $unsigned(_T_8715); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28779.4]
  assign _T_8717 = _T_8716[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28780.4]
  assign _T_8718 = _T_8712 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28782.4]
  assign _T_8720 = _T_8718 | _T_8704; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28784.4]
  assign _T_8722 = _T_8720 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28786.4]
  assign _T_8723 = _T_8722 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28787.4]
  assign _T_8724 = _T_8709 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28792.4]
  assign _T_8725 = _T_8704 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28793.4]
  assign _T_8726 = _T_8724 | _T_8725; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28794.4]
  assign _T_8728 = _T_8726 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28796.4]
  assign _T_8729 = _T_8728 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28797.4]
  assign _T_8740 = _T_2607 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28814.4]
  assign _T_8741 = _T_2867 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28815.4]
  assign _T_8743 = _T_8741 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28817.4]
  assign _T_8745 = _T_8735 + _T_8740; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28819.4]
  assign _T_8746 = _T_8745 - _T_8743; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28820.4]
  assign _T_8747 = $unsigned(_T_8746); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28821.4]
  assign _T_8748 = _T_8747[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28822.4]
  assign _T_8749 = _T_8743 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28824.4]
  assign _T_8751 = _T_8749 | _T_8735; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28826.4]
  assign _T_8753 = _T_8751 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28828.4]
  assign _T_8754 = _T_8753 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28829.4]
  assign _T_8755 = _T_8740 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28834.4]
  assign _T_8756 = _T_8735 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28835.4]
  assign _T_8757 = _T_8755 | _T_8756; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28836.4]
  assign _T_8759 = _T_8757 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28838.4]
  assign _T_8760 = _T_8759 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28839.4]
  assign _T_8771 = _T_2608 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28856.4]
  assign _T_8772 = _T_2868 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28857.4]
  assign _T_8774 = _T_8772 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28859.4]
  assign _T_8776 = _T_8766 + _T_8771; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28861.4]
  assign _T_8777 = _T_8776 - _T_8774; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28862.4]
  assign _T_8778 = $unsigned(_T_8777); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28863.4]
  assign _T_8779 = _T_8778[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28864.4]
  assign _T_8780 = _T_8774 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28866.4]
  assign _T_8782 = _T_8780 | _T_8766; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28868.4]
  assign _T_8784 = _T_8782 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28870.4]
  assign _T_8785 = _T_8784 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28871.4]
  assign _T_8786 = _T_8771 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28876.4]
  assign _T_8787 = _T_8766 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28877.4]
  assign _T_8788 = _T_8786 | _T_8787; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28878.4]
  assign _T_8790 = _T_8788 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28880.4]
  assign _T_8791 = _T_8790 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28881.4]
  assign _T_8802 = _T_2609 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28898.4]
  assign _T_8803 = _T_2869 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28899.4]
  assign _T_8805 = _T_8803 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28901.4]
  assign _T_8807 = _T_8797 + _T_8802; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28903.4]
  assign _T_8808 = _T_8807 - _T_8805; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28904.4]
  assign _T_8809 = $unsigned(_T_8808); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28905.4]
  assign _T_8810 = _T_8809[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28906.4]
  assign _T_8811 = _T_8805 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28908.4]
  assign _T_8813 = _T_8811 | _T_8797; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28910.4]
  assign _T_8815 = _T_8813 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28912.4]
  assign _T_8816 = _T_8815 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28913.4]
  assign _T_8817 = _T_8802 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28918.4]
  assign _T_8818 = _T_8797 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28919.4]
  assign _T_8819 = _T_8817 | _T_8818; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28920.4]
  assign _T_8821 = _T_8819 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28922.4]
  assign _T_8822 = _T_8821 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28923.4]
  assign _T_8833 = _T_2610 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28940.4]
  assign _T_8834 = _T_2870 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28941.4]
  assign _T_8836 = _T_8834 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28943.4]
  assign _T_8838 = _T_8828 + _T_8833; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28945.4]
  assign _T_8839 = _T_8838 - _T_8836; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28946.4]
  assign _T_8840 = $unsigned(_T_8839); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28947.4]
  assign _T_8841 = _T_8840[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28948.4]
  assign _T_8842 = _T_8836 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28950.4]
  assign _T_8844 = _T_8842 | _T_8828; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28952.4]
  assign _T_8846 = _T_8844 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28954.4]
  assign _T_8847 = _T_8846 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28955.4]
  assign _T_8848 = _T_8833 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@28960.4]
  assign _T_8849 = _T_8828 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@28961.4]
  assign _T_8850 = _T_8848 | _T_8849; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@28962.4]
  assign _T_8852 = _T_8850 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28964.4]
  assign _T_8853 = _T_8852 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28965.4]
  assign _T_8864 = _T_2611 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@28982.4]
  assign _T_8865 = _T_2871 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@28983.4]
  assign _T_8867 = _T_8865 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@28985.4]
  assign _T_8869 = _T_8859 + _T_8864; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@28987.4]
  assign _T_8870 = _T_8869 - _T_8867; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28988.4]
  assign _T_8871 = $unsigned(_T_8870); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28989.4]
  assign _T_8872 = _T_8871[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@28990.4]
  assign _T_8873 = _T_8867 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@28992.4]
  assign _T_8875 = _T_8873 | _T_8859; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@28994.4]
  assign _T_8877 = _T_8875 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28996.4]
  assign _T_8878 = _T_8877 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28997.4]
  assign _T_8879 = _T_8864 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29002.4]
  assign _T_8880 = _T_8859 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29003.4]
  assign _T_8881 = _T_8879 | _T_8880; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29004.4]
  assign _T_8883 = _T_8881 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29006.4]
  assign _T_8884 = _T_8883 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29007.4]
  assign _T_8895 = _T_2612 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29024.4]
  assign _T_8896 = _T_2872 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29025.4]
  assign _T_8898 = _T_8896 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29027.4]
  assign _T_8900 = _T_8890 + _T_8895; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29029.4]
  assign _T_8901 = _T_8900 - _T_8898; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29030.4]
  assign _T_8902 = $unsigned(_T_8901); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29031.4]
  assign _T_8903 = _T_8902[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29032.4]
  assign _T_8904 = _T_8898 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29034.4]
  assign _T_8906 = _T_8904 | _T_8890; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29036.4]
  assign _T_8908 = _T_8906 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29038.4]
  assign _T_8909 = _T_8908 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29039.4]
  assign _T_8910 = _T_8895 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29044.4]
  assign _T_8911 = _T_8890 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29045.4]
  assign _T_8912 = _T_8910 | _T_8911; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29046.4]
  assign _T_8914 = _T_8912 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29048.4]
  assign _T_8915 = _T_8914 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29049.4]
  assign _T_8926 = _T_2613 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29066.4]
  assign _T_8927 = _T_2873 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29067.4]
  assign _T_8929 = _T_8927 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29069.4]
  assign _T_8931 = _T_8921 + _T_8926; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29071.4]
  assign _T_8932 = _T_8931 - _T_8929; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29072.4]
  assign _T_8933 = $unsigned(_T_8932); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29073.4]
  assign _T_8934 = _T_8933[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29074.4]
  assign _T_8935 = _T_8929 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29076.4]
  assign _T_8937 = _T_8935 | _T_8921; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29078.4]
  assign _T_8939 = _T_8937 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29080.4]
  assign _T_8940 = _T_8939 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29081.4]
  assign _T_8941 = _T_8926 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29086.4]
  assign _T_8942 = _T_8921 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29087.4]
  assign _T_8943 = _T_8941 | _T_8942; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29088.4]
  assign _T_8945 = _T_8943 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29090.4]
  assign _T_8946 = _T_8945 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29091.4]
  assign _T_8957 = _T_2614 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29108.4]
  assign _T_8958 = _T_2874 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29109.4]
  assign _T_8960 = _T_8958 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29111.4]
  assign _T_8962 = _T_8952 + _T_8957; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29113.4]
  assign _T_8963 = _T_8962 - _T_8960; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29114.4]
  assign _T_8964 = $unsigned(_T_8963); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29115.4]
  assign _T_8965 = _T_8964[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29116.4]
  assign _T_8966 = _T_8960 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29118.4]
  assign _T_8968 = _T_8966 | _T_8952; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29120.4]
  assign _T_8970 = _T_8968 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29122.4]
  assign _T_8971 = _T_8970 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29123.4]
  assign _T_8972 = _T_8957 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29128.4]
  assign _T_8973 = _T_8952 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29129.4]
  assign _T_8974 = _T_8972 | _T_8973; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29130.4]
  assign _T_8976 = _T_8974 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29132.4]
  assign _T_8977 = _T_8976 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29133.4]
  assign _T_8988 = _T_2615 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29150.4]
  assign _T_8989 = _T_2875 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29151.4]
  assign _T_8991 = _T_8989 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29153.4]
  assign _T_8993 = _T_8983 + _T_8988; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29155.4]
  assign _T_8994 = _T_8993 - _T_8991; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29156.4]
  assign _T_8995 = $unsigned(_T_8994); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29157.4]
  assign _T_8996 = _T_8995[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29158.4]
  assign _T_8997 = _T_8991 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29160.4]
  assign _T_8999 = _T_8997 | _T_8983; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29162.4]
  assign _T_9001 = _T_8999 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29164.4]
  assign _T_9002 = _T_9001 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29165.4]
  assign _T_9003 = _T_8988 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29170.4]
  assign _T_9004 = _T_8983 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29171.4]
  assign _T_9005 = _T_9003 | _T_9004; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29172.4]
  assign _T_9007 = _T_9005 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29174.4]
  assign _T_9008 = _T_9007 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29175.4]
  assign _T_9019 = _T_2616 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29192.4]
  assign _T_9020 = _T_2876 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29193.4]
  assign _T_9022 = _T_9020 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29195.4]
  assign _T_9024 = _T_9014 + _T_9019; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29197.4]
  assign _T_9025 = _T_9024 - _T_9022; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29198.4]
  assign _T_9026 = $unsigned(_T_9025); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29199.4]
  assign _T_9027 = _T_9026[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29200.4]
  assign _T_9028 = _T_9022 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29202.4]
  assign _T_9030 = _T_9028 | _T_9014; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29204.4]
  assign _T_9032 = _T_9030 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29206.4]
  assign _T_9033 = _T_9032 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29207.4]
  assign _T_9034 = _T_9019 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29212.4]
  assign _T_9035 = _T_9014 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29213.4]
  assign _T_9036 = _T_9034 | _T_9035; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29214.4]
  assign _T_9038 = _T_9036 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29216.4]
  assign _T_9039 = _T_9038 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29217.4]
  assign _T_9050 = _T_2617 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29234.4]
  assign _T_9051 = _T_2877 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29235.4]
  assign _T_9053 = _T_9051 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29237.4]
  assign _T_9055 = _T_9045 + _T_9050; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29239.4]
  assign _T_9056 = _T_9055 - _T_9053; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29240.4]
  assign _T_9057 = $unsigned(_T_9056); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29241.4]
  assign _T_9058 = _T_9057[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29242.4]
  assign _T_9059 = _T_9053 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29244.4]
  assign _T_9061 = _T_9059 | _T_9045; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29246.4]
  assign _T_9063 = _T_9061 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29248.4]
  assign _T_9064 = _T_9063 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29249.4]
  assign _T_9065 = _T_9050 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29254.4]
  assign _T_9066 = _T_9045 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29255.4]
  assign _T_9067 = _T_9065 | _T_9066; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29256.4]
  assign _T_9069 = _T_9067 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29258.4]
  assign _T_9070 = _T_9069 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29259.4]
  assign _T_9081 = _T_2618 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29276.4]
  assign _T_9082 = _T_2878 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29277.4]
  assign _T_9084 = _T_9082 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29279.4]
  assign _T_9086 = _T_9076 + _T_9081; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29281.4]
  assign _T_9087 = _T_9086 - _T_9084; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29282.4]
  assign _T_9088 = $unsigned(_T_9087); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29283.4]
  assign _T_9089 = _T_9088[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29284.4]
  assign _T_9090 = _T_9084 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29286.4]
  assign _T_9092 = _T_9090 | _T_9076; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29288.4]
  assign _T_9094 = _T_9092 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29290.4]
  assign _T_9095 = _T_9094 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29291.4]
  assign _T_9096 = _T_9081 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29296.4]
  assign _T_9097 = _T_9076 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29297.4]
  assign _T_9098 = _T_9096 | _T_9097; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29298.4]
  assign _T_9100 = _T_9098 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29300.4]
  assign _T_9101 = _T_9100 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29301.4]
  assign _T_9112 = _T_2619 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29318.4]
  assign _T_9113 = _T_2879 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29319.4]
  assign _T_9115 = _T_9113 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29321.4]
  assign _T_9117 = _T_9107 + _T_9112; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29323.4]
  assign _T_9118 = _T_9117 - _T_9115; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29324.4]
  assign _T_9119 = $unsigned(_T_9118); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29325.4]
  assign _T_9120 = _T_9119[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29326.4]
  assign _T_9121 = _T_9115 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29328.4]
  assign _T_9123 = _T_9121 | _T_9107; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29330.4]
  assign _T_9125 = _T_9123 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29332.4]
  assign _T_9126 = _T_9125 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29333.4]
  assign _T_9127 = _T_9112 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29338.4]
  assign _T_9128 = _T_9107 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29339.4]
  assign _T_9129 = _T_9127 | _T_9128; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29340.4]
  assign _T_9131 = _T_9129 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29342.4]
  assign _T_9132 = _T_9131 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29343.4]
  assign _T_9143 = _T_2620 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29360.4]
  assign _T_9144 = _T_2880 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29361.4]
  assign _T_9146 = _T_9144 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29363.4]
  assign _T_9148 = _T_9138 + _T_9143; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29365.4]
  assign _T_9149 = _T_9148 - _T_9146; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29366.4]
  assign _T_9150 = $unsigned(_T_9149); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29367.4]
  assign _T_9151 = _T_9150[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29368.4]
  assign _T_9152 = _T_9146 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29370.4]
  assign _T_9154 = _T_9152 | _T_9138; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29372.4]
  assign _T_9156 = _T_9154 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29374.4]
  assign _T_9157 = _T_9156 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29375.4]
  assign _T_9158 = _T_9143 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29380.4]
  assign _T_9159 = _T_9138 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29381.4]
  assign _T_9160 = _T_9158 | _T_9159; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29382.4]
  assign _T_9162 = _T_9160 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29384.4]
  assign _T_9163 = _T_9162 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29385.4]
  assign _T_9174 = _T_2621 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29402.4]
  assign _T_9175 = _T_2881 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29403.4]
  assign _T_9177 = _T_9175 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29405.4]
  assign _T_9179 = _T_9169 + _T_9174; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29407.4]
  assign _T_9180 = _T_9179 - _T_9177; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29408.4]
  assign _T_9181 = $unsigned(_T_9180); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29409.4]
  assign _T_9182 = _T_9181[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29410.4]
  assign _T_9183 = _T_9177 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29412.4]
  assign _T_9185 = _T_9183 | _T_9169; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29414.4]
  assign _T_9187 = _T_9185 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29416.4]
  assign _T_9188 = _T_9187 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29417.4]
  assign _T_9189 = _T_9174 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29422.4]
  assign _T_9190 = _T_9169 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29423.4]
  assign _T_9191 = _T_9189 | _T_9190; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29424.4]
  assign _T_9193 = _T_9191 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29426.4]
  assign _T_9194 = _T_9193 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29427.4]
  assign _T_9205 = _T_2622 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29444.4]
  assign _T_9206 = _T_2882 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29445.4]
  assign _T_9208 = _T_9206 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29447.4]
  assign _T_9210 = _T_9200 + _T_9205; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29449.4]
  assign _T_9211 = _T_9210 - _T_9208; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29450.4]
  assign _T_9212 = $unsigned(_T_9211); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29451.4]
  assign _T_9213 = _T_9212[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29452.4]
  assign _T_9214 = _T_9208 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29454.4]
  assign _T_9216 = _T_9214 | _T_9200; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29456.4]
  assign _T_9218 = _T_9216 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29458.4]
  assign _T_9219 = _T_9218 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29459.4]
  assign _T_9220 = _T_9205 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29464.4]
  assign _T_9221 = _T_9200 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29465.4]
  assign _T_9222 = _T_9220 | _T_9221; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29466.4]
  assign _T_9224 = _T_9222 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29468.4]
  assign _T_9225 = _T_9224 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29469.4]
  assign _T_9236 = _T_2623 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29486.4]
  assign _T_9237 = _T_2883 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29487.4]
  assign _T_9239 = _T_9237 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29489.4]
  assign _T_9241 = _T_9231 + _T_9236; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29491.4]
  assign _T_9242 = _T_9241 - _T_9239; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29492.4]
  assign _T_9243 = $unsigned(_T_9242); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29493.4]
  assign _T_9244 = _T_9243[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29494.4]
  assign _T_9245 = _T_9239 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29496.4]
  assign _T_9247 = _T_9245 | _T_9231; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29498.4]
  assign _T_9249 = _T_9247 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29500.4]
  assign _T_9250 = _T_9249 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29501.4]
  assign _T_9251 = _T_9236 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29506.4]
  assign _T_9252 = _T_9231 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29507.4]
  assign _T_9253 = _T_9251 | _T_9252; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29508.4]
  assign _T_9255 = _T_9253 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29510.4]
  assign _T_9256 = _T_9255 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29511.4]
  assign _T_9267 = _T_2624 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29528.4]
  assign _T_9268 = _T_2884 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29529.4]
  assign _T_9270 = _T_9268 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29531.4]
  assign _T_9272 = _T_9262 + _T_9267; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29533.4]
  assign _T_9273 = _T_9272 - _T_9270; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29534.4]
  assign _T_9274 = $unsigned(_T_9273); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29535.4]
  assign _T_9275 = _T_9274[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29536.4]
  assign _T_9276 = _T_9270 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29538.4]
  assign _T_9278 = _T_9276 | _T_9262; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29540.4]
  assign _T_9280 = _T_9278 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29542.4]
  assign _T_9281 = _T_9280 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29543.4]
  assign _T_9282 = _T_9267 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29548.4]
  assign _T_9283 = _T_9262 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29549.4]
  assign _T_9284 = _T_9282 | _T_9283; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29550.4]
  assign _T_9286 = _T_9284 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29552.4]
  assign _T_9287 = _T_9286 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29553.4]
  assign _T_9298 = _T_2625 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29570.4]
  assign _T_9299 = _T_2885 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29571.4]
  assign _T_9301 = _T_9299 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29573.4]
  assign _T_9303 = _T_9293 + _T_9298; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29575.4]
  assign _T_9304 = _T_9303 - _T_9301; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29576.4]
  assign _T_9305 = $unsigned(_T_9304); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29577.4]
  assign _T_9306 = _T_9305[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29578.4]
  assign _T_9307 = _T_9301 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29580.4]
  assign _T_9309 = _T_9307 | _T_9293; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29582.4]
  assign _T_9311 = _T_9309 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29584.4]
  assign _T_9312 = _T_9311 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29585.4]
  assign _T_9313 = _T_9298 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29590.4]
  assign _T_9314 = _T_9293 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29591.4]
  assign _T_9315 = _T_9313 | _T_9314; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29592.4]
  assign _T_9317 = _T_9315 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29594.4]
  assign _T_9318 = _T_9317 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29595.4]
  assign _T_9329 = _T_2626 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29612.4]
  assign _T_9330 = _T_2886 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29613.4]
  assign _T_9332 = _T_9330 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29615.4]
  assign _T_9334 = _T_9324 + _T_9329; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29617.4]
  assign _T_9335 = _T_9334 - _T_9332; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29618.4]
  assign _T_9336 = $unsigned(_T_9335); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29619.4]
  assign _T_9337 = _T_9336[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29620.4]
  assign _T_9338 = _T_9332 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29622.4]
  assign _T_9340 = _T_9338 | _T_9324; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29624.4]
  assign _T_9342 = _T_9340 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29626.4]
  assign _T_9343 = _T_9342 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29627.4]
  assign _T_9344 = _T_9329 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29632.4]
  assign _T_9345 = _T_9324 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29633.4]
  assign _T_9346 = _T_9344 | _T_9345; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29634.4]
  assign _T_9348 = _T_9346 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29636.4]
  assign _T_9349 = _T_9348 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29637.4]
  assign _T_9360 = _T_2627 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29654.4]
  assign _T_9361 = _T_2887 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29655.4]
  assign _T_9363 = _T_9361 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29657.4]
  assign _T_9365 = _T_9355 + _T_9360; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29659.4]
  assign _T_9366 = _T_9365 - _T_9363; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29660.4]
  assign _T_9367 = $unsigned(_T_9366); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29661.4]
  assign _T_9368 = _T_9367[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29662.4]
  assign _T_9369 = _T_9363 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29664.4]
  assign _T_9371 = _T_9369 | _T_9355; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29666.4]
  assign _T_9373 = _T_9371 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29668.4]
  assign _T_9374 = _T_9373 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29669.4]
  assign _T_9375 = _T_9360 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29674.4]
  assign _T_9376 = _T_9355 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29675.4]
  assign _T_9377 = _T_9375 | _T_9376; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29676.4]
  assign _T_9379 = _T_9377 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29678.4]
  assign _T_9380 = _T_9379 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29679.4]
  assign _T_9391 = _T_2628 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29696.4]
  assign _T_9392 = _T_2888 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29697.4]
  assign _T_9394 = _T_9392 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29699.4]
  assign _T_9396 = _T_9386 + _T_9391; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29701.4]
  assign _T_9397 = _T_9396 - _T_9394; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29702.4]
  assign _T_9398 = $unsigned(_T_9397); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29703.4]
  assign _T_9399 = _T_9398[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29704.4]
  assign _T_9400 = _T_9394 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29706.4]
  assign _T_9402 = _T_9400 | _T_9386; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29708.4]
  assign _T_9404 = _T_9402 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29710.4]
  assign _T_9405 = _T_9404 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29711.4]
  assign _T_9406 = _T_9391 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29716.4]
  assign _T_9407 = _T_9386 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29717.4]
  assign _T_9408 = _T_9406 | _T_9407; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29718.4]
  assign _T_9410 = _T_9408 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29720.4]
  assign _T_9411 = _T_9410 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29721.4]
  assign _T_9422 = _T_2629 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29738.4]
  assign _T_9423 = _T_2889 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29739.4]
  assign _T_9425 = _T_9423 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29741.4]
  assign _T_9427 = _T_9417 + _T_9422; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29743.4]
  assign _T_9428 = _T_9427 - _T_9425; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29744.4]
  assign _T_9429 = $unsigned(_T_9428); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29745.4]
  assign _T_9430 = _T_9429[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29746.4]
  assign _T_9431 = _T_9425 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29748.4]
  assign _T_9433 = _T_9431 | _T_9417; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29750.4]
  assign _T_9435 = _T_9433 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29752.4]
  assign _T_9436 = _T_9435 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29753.4]
  assign _T_9437 = _T_9422 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29758.4]
  assign _T_9438 = _T_9417 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29759.4]
  assign _T_9439 = _T_9437 | _T_9438; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29760.4]
  assign _T_9441 = _T_9439 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29762.4]
  assign _T_9442 = _T_9441 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29763.4]
  assign _T_9453 = _T_2630 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29780.4]
  assign _T_9454 = _T_2890 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29781.4]
  assign _T_9456 = _T_9454 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29783.4]
  assign _T_9458 = _T_9448 + _T_9453; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29785.4]
  assign _T_9459 = _T_9458 - _T_9456; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29786.4]
  assign _T_9460 = $unsigned(_T_9459); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29787.4]
  assign _T_9461 = _T_9460[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29788.4]
  assign _T_9462 = _T_9456 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29790.4]
  assign _T_9464 = _T_9462 | _T_9448; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29792.4]
  assign _T_9466 = _T_9464 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29794.4]
  assign _T_9467 = _T_9466 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29795.4]
  assign _T_9468 = _T_9453 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29800.4]
  assign _T_9469 = _T_9448 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29801.4]
  assign _T_9470 = _T_9468 | _T_9469; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29802.4]
  assign _T_9472 = _T_9470 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29804.4]
  assign _T_9473 = _T_9472 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29805.4]
  assign _T_9484 = _T_2631 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29822.4]
  assign _T_9485 = _T_2891 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29823.4]
  assign _T_9487 = _T_9485 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29825.4]
  assign _T_9489 = _T_9479 + _T_9484; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29827.4]
  assign _T_9490 = _T_9489 - _T_9487; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29828.4]
  assign _T_9491 = $unsigned(_T_9490); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29829.4]
  assign _T_9492 = _T_9491[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29830.4]
  assign _T_9493 = _T_9487 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29832.4]
  assign _T_9495 = _T_9493 | _T_9479; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29834.4]
  assign _T_9497 = _T_9495 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29836.4]
  assign _T_9498 = _T_9497 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29837.4]
  assign _T_9499 = _T_9484 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29842.4]
  assign _T_9500 = _T_9479 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29843.4]
  assign _T_9501 = _T_9499 | _T_9500; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29844.4]
  assign _T_9503 = _T_9501 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29846.4]
  assign _T_9504 = _T_9503 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29847.4]
  assign _T_9515 = _T_2632 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29864.4]
  assign _T_9516 = _T_2892 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29865.4]
  assign _T_9518 = _T_9516 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29867.4]
  assign _T_9520 = _T_9510 + _T_9515; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29869.4]
  assign _T_9521 = _T_9520 - _T_9518; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29870.4]
  assign _T_9522 = $unsigned(_T_9521); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29871.4]
  assign _T_9523 = _T_9522[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29872.4]
  assign _T_9524 = _T_9518 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29874.4]
  assign _T_9526 = _T_9524 | _T_9510; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29876.4]
  assign _T_9528 = _T_9526 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29878.4]
  assign _T_9529 = _T_9528 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29879.4]
  assign _T_9530 = _T_9515 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29884.4]
  assign _T_9531 = _T_9510 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29885.4]
  assign _T_9532 = _T_9530 | _T_9531; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29886.4]
  assign _T_9534 = _T_9532 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29888.4]
  assign _T_9535 = _T_9534 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29889.4]
  assign _T_9546 = _T_2633 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29906.4]
  assign _T_9547 = _T_2893 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29907.4]
  assign _T_9549 = _T_9547 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29909.4]
  assign _T_9551 = _T_9541 + _T_9546; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29911.4]
  assign _T_9552 = _T_9551 - _T_9549; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29912.4]
  assign _T_9553 = $unsigned(_T_9552); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29913.4]
  assign _T_9554 = _T_9553[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29914.4]
  assign _T_9555 = _T_9549 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29916.4]
  assign _T_9557 = _T_9555 | _T_9541; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29918.4]
  assign _T_9559 = _T_9557 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29920.4]
  assign _T_9560 = _T_9559 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29921.4]
  assign _T_9561 = _T_9546 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29926.4]
  assign _T_9562 = _T_9541 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29927.4]
  assign _T_9563 = _T_9561 | _T_9562; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29928.4]
  assign _T_9565 = _T_9563 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29930.4]
  assign _T_9566 = _T_9565 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29931.4]
  assign _T_9577 = _T_2634 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29948.4]
  assign _T_9578 = _T_2894 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29949.4]
  assign _T_9580 = _T_9578 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29951.4]
  assign _T_9582 = _T_9572 + _T_9577; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29953.4]
  assign _T_9583 = _T_9582 - _T_9580; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29954.4]
  assign _T_9584 = $unsigned(_T_9583); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29955.4]
  assign _T_9585 = _T_9584[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29956.4]
  assign _T_9586 = _T_9580 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@29958.4]
  assign _T_9588 = _T_9586 | _T_9572; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@29960.4]
  assign _T_9590 = _T_9588 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29962.4]
  assign _T_9591 = _T_9590 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29963.4]
  assign _T_9592 = _T_9577 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@29968.4]
  assign _T_9593 = _T_9572 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@29969.4]
  assign _T_9594 = _T_9592 | _T_9593; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@29970.4]
  assign _T_9596 = _T_9594 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29972.4]
  assign _T_9597 = _T_9596 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29973.4]
  assign _T_9608 = _T_2635 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@29990.4]
  assign _T_9609 = _T_2895 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@29991.4]
  assign _T_9611 = _T_9609 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@29993.4]
  assign _T_9613 = _T_9603 + _T_9608; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@29995.4]
  assign _T_9614 = _T_9613 - _T_9611; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29996.4]
  assign _T_9615 = $unsigned(_T_9614); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29997.4]
  assign _T_9616 = _T_9615[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@29998.4]
  assign _T_9617 = _T_9611 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30000.4]
  assign _T_9619 = _T_9617 | _T_9603; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30002.4]
  assign _T_9621 = _T_9619 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30004.4]
  assign _T_9622 = _T_9621 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30005.4]
  assign _T_9623 = _T_9608 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30010.4]
  assign _T_9624 = _T_9603 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30011.4]
  assign _T_9625 = _T_9623 | _T_9624; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30012.4]
  assign _T_9627 = _T_9625 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30014.4]
  assign _T_9628 = _T_9627 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30015.4]
  assign _T_9639 = _T_2636 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30032.4]
  assign _T_9640 = _T_2896 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30033.4]
  assign _T_9642 = _T_9640 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30035.4]
  assign _T_9644 = _T_9634 + _T_9639; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30037.4]
  assign _T_9645 = _T_9644 - _T_9642; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30038.4]
  assign _T_9646 = $unsigned(_T_9645); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30039.4]
  assign _T_9647 = _T_9646[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30040.4]
  assign _T_9648 = _T_9642 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30042.4]
  assign _T_9650 = _T_9648 | _T_9634; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30044.4]
  assign _T_9652 = _T_9650 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30046.4]
  assign _T_9653 = _T_9652 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30047.4]
  assign _T_9654 = _T_9639 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30052.4]
  assign _T_9655 = _T_9634 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30053.4]
  assign _T_9656 = _T_9654 | _T_9655; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30054.4]
  assign _T_9658 = _T_9656 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30056.4]
  assign _T_9659 = _T_9658 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30057.4]
  assign _T_9670 = _T_2637 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30074.4]
  assign _T_9671 = _T_2897 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30075.4]
  assign _T_9673 = _T_9671 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30077.4]
  assign _T_9675 = _T_9665 + _T_9670; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30079.4]
  assign _T_9676 = _T_9675 - _T_9673; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30080.4]
  assign _T_9677 = $unsigned(_T_9676); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30081.4]
  assign _T_9678 = _T_9677[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30082.4]
  assign _T_9679 = _T_9673 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30084.4]
  assign _T_9681 = _T_9679 | _T_9665; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30086.4]
  assign _T_9683 = _T_9681 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30088.4]
  assign _T_9684 = _T_9683 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30089.4]
  assign _T_9685 = _T_9670 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30094.4]
  assign _T_9686 = _T_9665 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30095.4]
  assign _T_9687 = _T_9685 | _T_9686; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30096.4]
  assign _T_9689 = _T_9687 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30098.4]
  assign _T_9690 = _T_9689 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30099.4]
  assign _T_9701 = _T_2638 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30116.4]
  assign _T_9702 = _T_2898 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30117.4]
  assign _T_9704 = _T_9702 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30119.4]
  assign _T_9706 = _T_9696 + _T_9701; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30121.4]
  assign _T_9707 = _T_9706 - _T_9704; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30122.4]
  assign _T_9708 = $unsigned(_T_9707); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30123.4]
  assign _T_9709 = _T_9708[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30124.4]
  assign _T_9710 = _T_9704 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30126.4]
  assign _T_9712 = _T_9710 | _T_9696; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30128.4]
  assign _T_9714 = _T_9712 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30130.4]
  assign _T_9715 = _T_9714 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30131.4]
  assign _T_9716 = _T_9701 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30136.4]
  assign _T_9717 = _T_9696 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30137.4]
  assign _T_9718 = _T_9716 | _T_9717; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30138.4]
  assign _T_9720 = _T_9718 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30140.4]
  assign _T_9721 = _T_9720 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30141.4]
  assign _T_9732 = _T_2639 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30158.4]
  assign _T_9733 = _T_2899 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30159.4]
  assign _T_9735 = _T_9733 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30161.4]
  assign _T_9737 = _T_9727 + _T_9732; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30163.4]
  assign _T_9738 = _T_9737 - _T_9735; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30164.4]
  assign _T_9739 = $unsigned(_T_9738); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30165.4]
  assign _T_9740 = _T_9739[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30166.4]
  assign _T_9741 = _T_9735 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30168.4]
  assign _T_9743 = _T_9741 | _T_9727; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30170.4]
  assign _T_9745 = _T_9743 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30172.4]
  assign _T_9746 = _T_9745 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30173.4]
  assign _T_9747 = _T_9732 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30178.4]
  assign _T_9748 = _T_9727 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30179.4]
  assign _T_9749 = _T_9747 | _T_9748; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30180.4]
  assign _T_9751 = _T_9749 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30182.4]
  assign _T_9752 = _T_9751 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30183.4]
  assign _T_9763 = _T_2640 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30200.4]
  assign _T_9764 = _T_2900 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30201.4]
  assign _T_9766 = _T_9764 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30203.4]
  assign _T_9768 = _T_9758 + _T_9763; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30205.4]
  assign _T_9769 = _T_9768 - _T_9766; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30206.4]
  assign _T_9770 = $unsigned(_T_9769); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30207.4]
  assign _T_9771 = _T_9770[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30208.4]
  assign _T_9772 = _T_9766 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30210.4]
  assign _T_9774 = _T_9772 | _T_9758; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30212.4]
  assign _T_9776 = _T_9774 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30214.4]
  assign _T_9777 = _T_9776 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30215.4]
  assign _T_9778 = _T_9763 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30220.4]
  assign _T_9779 = _T_9758 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30221.4]
  assign _T_9780 = _T_9778 | _T_9779; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30222.4]
  assign _T_9782 = _T_9780 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30224.4]
  assign _T_9783 = _T_9782 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30225.4]
  assign _T_9794 = _T_2641 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30242.4]
  assign _T_9795 = _T_2901 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30243.4]
  assign _T_9797 = _T_9795 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30245.4]
  assign _T_9799 = _T_9789 + _T_9794; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30247.4]
  assign _T_9800 = _T_9799 - _T_9797; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30248.4]
  assign _T_9801 = $unsigned(_T_9800); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30249.4]
  assign _T_9802 = _T_9801[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30250.4]
  assign _T_9803 = _T_9797 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30252.4]
  assign _T_9805 = _T_9803 | _T_9789; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30254.4]
  assign _T_9807 = _T_9805 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30256.4]
  assign _T_9808 = _T_9807 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30257.4]
  assign _T_9809 = _T_9794 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30262.4]
  assign _T_9810 = _T_9789 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30263.4]
  assign _T_9811 = _T_9809 | _T_9810; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30264.4]
  assign _T_9813 = _T_9811 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30266.4]
  assign _T_9814 = _T_9813 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30267.4]
  assign _T_9825 = _T_2642 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30284.4]
  assign _T_9826 = _T_2902 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30285.4]
  assign _T_9828 = _T_9826 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30287.4]
  assign _T_9830 = _T_9820 + _T_9825; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30289.4]
  assign _T_9831 = _T_9830 - _T_9828; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30290.4]
  assign _T_9832 = $unsigned(_T_9831); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30291.4]
  assign _T_9833 = _T_9832[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30292.4]
  assign _T_9834 = _T_9828 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30294.4]
  assign _T_9836 = _T_9834 | _T_9820; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30296.4]
  assign _T_9838 = _T_9836 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30298.4]
  assign _T_9839 = _T_9838 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30299.4]
  assign _T_9840 = _T_9825 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30304.4]
  assign _T_9841 = _T_9820 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30305.4]
  assign _T_9842 = _T_9840 | _T_9841; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30306.4]
  assign _T_9844 = _T_9842 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30308.4]
  assign _T_9845 = _T_9844 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30309.4]
  assign _T_9856 = _T_2643 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30326.4]
  assign _T_9857 = _T_2903 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30327.4]
  assign _T_9859 = _T_9857 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30329.4]
  assign _T_9861 = _T_9851 + _T_9856; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30331.4]
  assign _T_9862 = _T_9861 - _T_9859; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30332.4]
  assign _T_9863 = $unsigned(_T_9862); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30333.4]
  assign _T_9864 = _T_9863[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30334.4]
  assign _T_9865 = _T_9859 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30336.4]
  assign _T_9867 = _T_9865 | _T_9851; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30338.4]
  assign _T_9869 = _T_9867 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30340.4]
  assign _T_9870 = _T_9869 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30341.4]
  assign _T_9871 = _T_9856 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30346.4]
  assign _T_9872 = _T_9851 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30347.4]
  assign _T_9873 = _T_9871 | _T_9872; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30348.4]
  assign _T_9875 = _T_9873 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30350.4]
  assign _T_9876 = _T_9875 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30351.4]
  assign _T_9887 = _T_2644 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30368.4]
  assign _T_9888 = _T_2904 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30369.4]
  assign _T_9890 = _T_9888 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30371.4]
  assign _T_9892 = _T_9882 + _T_9887; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30373.4]
  assign _T_9893 = _T_9892 - _T_9890; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30374.4]
  assign _T_9894 = $unsigned(_T_9893); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30375.4]
  assign _T_9895 = _T_9894[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30376.4]
  assign _T_9896 = _T_9890 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30378.4]
  assign _T_9898 = _T_9896 | _T_9882; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30380.4]
  assign _T_9900 = _T_9898 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30382.4]
  assign _T_9901 = _T_9900 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30383.4]
  assign _T_9902 = _T_9887 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30388.4]
  assign _T_9903 = _T_9882 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30389.4]
  assign _T_9904 = _T_9902 | _T_9903; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30390.4]
  assign _T_9906 = _T_9904 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30392.4]
  assign _T_9907 = _T_9906 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30393.4]
  assign _T_9918 = _T_2645 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30410.4]
  assign _T_9919 = _T_2905 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30411.4]
  assign _T_9921 = _T_9919 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30413.4]
  assign _T_9923 = _T_9913 + _T_9918; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30415.4]
  assign _T_9924 = _T_9923 - _T_9921; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30416.4]
  assign _T_9925 = $unsigned(_T_9924); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30417.4]
  assign _T_9926 = _T_9925[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30418.4]
  assign _T_9927 = _T_9921 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30420.4]
  assign _T_9929 = _T_9927 | _T_9913; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30422.4]
  assign _T_9931 = _T_9929 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30424.4]
  assign _T_9932 = _T_9931 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30425.4]
  assign _T_9933 = _T_9918 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30430.4]
  assign _T_9934 = _T_9913 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30431.4]
  assign _T_9935 = _T_9933 | _T_9934; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30432.4]
  assign _T_9937 = _T_9935 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30434.4]
  assign _T_9938 = _T_9937 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30435.4]
  assign _T_9949 = _T_2646 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30452.4]
  assign _T_9950 = _T_2906 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30453.4]
  assign _T_9952 = _T_9950 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30455.4]
  assign _T_9954 = _T_9944 + _T_9949; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30457.4]
  assign _T_9955 = _T_9954 - _T_9952; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30458.4]
  assign _T_9956 = $unsigned(_T_9955); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30459.4]
  assign _T_9957 = _T_9956[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30460.4]
  assign _T_9958 = _T_9952 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30462.4]
  assign _T_9960 = _T_9958 | _T_9944; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30464.4]
  assign _T_9962 = _T_9960 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30466.4]
  assign _T_9963 = _T_9962 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30467.4]
  assign _T_9964 = _T_9949 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30472.4]
  assign _T_9965 = _T_9944 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30473.4]
  assign _T_9966 = _T_9964 | _T_9965; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30474.4]
  assign _T_9968 = _T_9966 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30476.4]
  assign _T_9969 = _T_9968 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30477.4]
  assign _T_9980 = _T_2647 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30494.4]
  assign _T_9981 = _T_2907 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30495.4]
  assign _T_9983 = _T_9981 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30497.4]
  assign _T_9985 = _T_9975 + _T_9980; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30499.4]
  assign _T_9986 = _T_9985 - _T_9983; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30500.4]
  assign _T_9987 = $unsigned(_T_9986); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30501.4]
  assign _T_9988 = _T_9987[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30502.4]
  assign _T_9989 = _T_9983 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30504.4]
  assign _T_9991 = _T_9989 | _T_9975; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30506.4]
  assign _T_9993 = _T_9991 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30508.4]
  assign _T_9994 = _T_9993 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30509.4]
  assign _T_9995 = _T_9980 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30514.4]
  assign _T_9996 = _T_9975 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30515.4]
  assign _T_9997 = _T_9995 | _T_9996; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30516.4]
  assign _T_9999 = _T_9997 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30518.4]
  assign _T_10000 = _T_9999 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30519.4]
  assign _T_10011 = _T_2648 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30536.4]
  assign _T_10012 = _T_2908 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30537.4]
  assign _T_10014 = _T_10012 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30539.4]
  assign _T_10016 = _T_10006 + _T_10011; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30541.4]
  assign _T_10017 = _T_10016 - _T_10014; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30542.4]
  assign _T_10018 = $unsigned(_T_10017); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30543.4]
  assign _T_10019 = _T_10018[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30544.4]
  assign _T_10020 = _T_10014 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30546.4]
  assign _T_10022 = _T_10020 | _T_10006; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30548.4]
  assign _T_10024 = _T_10022 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30550.4]
  assign _T_10025 = _T_10024 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30551.4]
  assign _T_10026 = _T_10011 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30556.4]
  assign _T_10027 = _T_10006 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30557.4]
  assign _T_10028 = _T_10026 | _T_10027; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30558.4]
  assign _T_10030 = _T_10028 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30560.4]
  assign _T_10031 = _T_10030 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30561.4]
  assign _T_10042 = _T_2649 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30578.4]
  assign _T_10043 = _T_2909 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30579.4]
  assign _T_10045 = _T_10043 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30581.4]
  assign _T_10047 = _T_10037 + _T_10042; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30583.4]
  assign _T_10048 = _T_10047 - _T_10045; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30584.4]
  assign _T_10049 = $unsigned(_T_10048); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30585.4]
  assign _T_10050 = _T_10049[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30586.4]
  assign _T_10051 = _T_10045 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30588.4]
  assign _T_10053 = _T_10051 | _T_10037; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30590.4]
  assign _T_10055 = _T_10053 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30592.4]
  assign _T_10056 = _T_10055 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30593.4]
  assign _T_10057 = _T_10042 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30598.4]
  assign _T_10058 = _T_10037 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30599.4]
  assign _T_10059 = _T_10057 | _T_10058; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30600.4]
  assign _T_10061 = _T_10059 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30602.4]
  assign _T_10062 = _T_10061 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30603.4]
  assign _T_10073 = _T_2650 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30620.4]
  assign _T_10074 = _T_2910 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30621.4]
  assign _T_10076 = _T_10074 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30623.4]
  assign _T_10078 = _T_10068 + _T_10073; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30625.4]
  assign _T_10079 = _T_10078 - _T_10076; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30626.4]
  assign _T_10080 = $unsigned(_T_10079); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30627.4]
  assign _T_10081 = _T_10080[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30628.4]
  assign _T_10082 = _T_10076 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30630.4]
  assign _T_10084 = _T_10082 | _T_10068; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30632.4]
  assign _T_10086 = _T_10084 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30634.4]
  assign _T_10087 = _T_10086 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30635.4]
  assign _T_10088 = _T_10073 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30640.4]
  assign _T_10089 = _T_10068 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30641.4]
  assign _T_10090 = _T_10088 | _T_10089; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30642.4]
  assign _T_10092 = _T_10090 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30644.4]
  assign _T_10093 = _T_10092 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30645.4]
  assign _T_10104 = _T_2651 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30662.4]
  assign _T_10105 = _T_2911 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30663.4]
  assign _T_10107 = _T_10105 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30665.4]
  assign _T_10109 = _T_10099 + _T_10104; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30667.4]
  assign _T_10110 = _T_10109 - _T_10107; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30668.4]
  assign _T_10111 = $unsigned(_T_10110); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30669.4]
  assign _T_10112 = _T_10111[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30670.4]
  assign _T_10113 = _T_10107 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30672.4]
  assign _T_10115 = _T_10113 | _T_10099; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30674.4]
  assign _T_10117 = _T_10115 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30676.4]
  assign _T_10118 = _T_10117 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30677.4]
  assign _T_10119 = _T_10104 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30682.4]
  assign _T_10120 = _T_10099 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30683.4]
  assign _T_10121 = _T_10119 | _T_10120; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30684.4]
  assign _T_10123 = _T_10121 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30686.4]
  assign _T_10124 = _T_10123 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30687.4]
  assign _T_10135 = _T_2652 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30704.4]
  assign _T_10136 = _T_2912 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30705.4]
  assign _T_10138 = _T_10136 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30707.4]
  assign _T_10140 = _T_10130 + _T_10135; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30709.4]
  assign _T_10141 = _T_10140 - _T_10138; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30710.4]
  assign _T_10142 = $unsigned(_T_10141); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30711.4]
  assign _T_10143 = _T_10142[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30712.4]
  assign _T_10144 = _T_10138 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30714.4]
  assign _T_10146 = _T_10144 | _T_10130; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30716.4]
  assign _T_10148 = _T_10146 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30718.4]
  assign _T_10149 = _T_10148 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30719.4]
  assign _T_10150 = _T_10135 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30724.4]
  assign _T_10151 = _T_10130 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30725.4]
  assign _T_10152 = _T_10150 | _T_10151; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30726.4]
  assign _T_10154 = _T_10152 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30728.4]
  assign _T_10155 = _T_10154 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30729.4]
  assign _T_10166 = _T_2653 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30746.4]
  assign _T_10167 = _T_2913 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30747.4]
  assign _T_10169 = _T_10167 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30749.4]
  assign _T_10171 = _T_10161 + _T_10166; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30751.4]
  assign _T_10172 = _T_10171 - _T_10169; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30752.4]
  assign _T_10173 = $unsigned(_T_10172); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30753.4]
  assign _T_10174 = _T_10173[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30754.4]
  assign _T_10175 = _T_10169 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30756.4]
  assign _T_10177 = _T_10175 | _T_10161; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30758.4]
  assign _T_10179 = _T_10177 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30760.4]
  assign _T_10180 = _T_10179 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30761.4]
  assign _T_10181 = _T_10166 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30766.4]
  assign _T_10182 = _T_10161 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30767.4]
  assign _T_10183 = _T_10181 | _T_10182; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30768.4]
  assign _T_10185 = _T_10183 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30770.4]
  assign _T_10186 = _T_10185 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30771.4]
  assign _T_10197 = _T_2654 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30788.4]
  assign _T_10198 = _T_2914 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30789.4]
  assign _T_10200 = _T_10198 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30791.4]
  assign _T_10202 = _T_10192 + _T_10197; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30793.4]
  assign _T_10203 = _T_10202 - _T_10200; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30794.4]
  assign _T_10204 = $unsigned(_T_10203); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30795.4]
  assign _T_10205 = _T_10204[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30796.4]
  assign _T_10206 = _T_10200 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30798.4]
  assign _T_10208 = _T_10206 | _T_10192; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30800.4]
  assign _T_10210 = _T_10208 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30802.4]
  assign _T_10211 = _T_10210 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30803.4]
  assign _T_10212 = _T_10197 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30808.4]
  assign _T_10213 = _T_10192 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30809.4]
  assign _T_10214 = _T_10212 | _T_10213; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30810.4]
  assign _T_10216 = _T_10214 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30812.4]
  assign _T_10217 = _T_10216 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30813.4]
  assign _T_10228 = _T_2655 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30830.4]
  assign _T_10229 = _T_2915 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30831.4]
  assign _T_10231 = _T_10229 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30833.4]
  assign _T_10233 = _T_10223 + _T_10228; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30835.4]
  assign _T_10234 = _T_10233 - _T_10231; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30836.4]
  assign _T_10235 = $unsigned(_T_10234); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30837.4]
  assign _T_10236 = _T_10235[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30838.4]
  assign _T_10237 = _T_10231 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30840.4]
  assign _T_10239 = _T_10237 | _T_10223; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30842.4]
  assign _T_10241 = _T_10239 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30844.4]
  assign _T_10242 = _T_10241 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30845.4]
  assign _T_10243 = _T_10228 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30850.4]
  assign _T_10244 = _T_10223 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30851.4]
  assign _T_10245 = _T_10243 | _T_10244; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30852.4]
  assign _T_10247 = _T_10245 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30854.4]
  assign _T_10248 = _T_10247 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30855.4]
  assign _T_10259 = _T_2656 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30872.4]
  assign _T_10260 = _T_2916 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30873.4]
  assign _T_10262 = _T_10260 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30875.4]
  assign _T_10264 = _T_10254 + _T_10259; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30877.4]
  assign _T_10265 = _T_10264 - _T_10262; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30878.4]
  assign _T_10266 = $unsigned(_T_10265); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30879.4]
  assign _T_10267 = _T_10266[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30880.4]
  assign _T_10268 = _T_10262 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30882.4]
  assign _T_10270 = _T_10268 | _T_10254; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30884.4]
  assign _T_10272 = _T_10270 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30886.4]
  assign _T_10273 = _T_10272 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30887.4]
  assign _T_10274 = _T_10259 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30892.4]
  assign _T_10275 = _T_10254 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30893.4]
  assign _T_10276 = _T_10274 | _T_10275; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30894.4]
  assign _T_10278 = _T_10276 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30896.4]
  assign _T_10279 = _T_10278 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30897.4]
  assign _T_10290 = _T_2657 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30914.4]
  assign _T_10291 = _T_2917 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30915.4]
  assign _T_10293 = _T_10291 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30917.4]
  assign _T_10295 = _T_10285 + _T_10290; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30919.4]
  assign _T_10296 = _T_10295 - _T_10293; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30920.4]
  assign _T_10297 = $unsigned(_T_10296); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30921.4]
  assign _T_10298 = _T_10297[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30922.4]
  assign _T_10299 = _T_10293 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30924.4]
  assign _T_10301 = _T_10299 | _T_10285; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30926.4]
  assign _T_10303 = _T_10301 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30928.4]
  assign _T_10304 = _T_10303 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30929.4]
  assign _T_10305 = _T_10290 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30934.4]
  assign _T_10306 = _T_10285 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30935.4]
  assign _T_10307 = _T_10305 | _T_10306; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30936.4]
  assign _T_10309 = _T_10307 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30938.4]
  assign _T_10310 = _T_10309 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30939.4]
  assign _T_10321 = _T_2658 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30956.4]
  assign _T_10322 = _T_2918 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30957.4]
  assign _T_10324 = _T_10322 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@30959.4]
  assign _T_10326 = _T_10316 + _T_10321; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@30961.4]
  assign _T_10327 = _T_10326 - _T_10324; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30962.4]
  assign _T_10328 = $unsigned(_T_10327); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30963.4]
  assign _T_10329 = _T_10328[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@30964.4]
  assign _T_10330 = _T_10324 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@30966.4]
  assign _T_10332 = _T_10330 | _T_10316; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@30968.4]
  assign _T_10334 = _T_10332 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30970.4]
  assign _T_10335 = _T_10334 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30971.4]
  assign _T_10336 = _T_10321 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@30976.4]
  assign _T_10337 = _T_10316 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@30977.4]
  assign _T_10338 = _T_10336 | _T_10337; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@30978.4]
  assign _T_10340 = _T_10338 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30980.4]
  assign _T_10341 = _T_10340 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30981.4]
  assign _T_10352 = _T_2659 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@30998.4]
  assign _T_10353 = _T_2919 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@30999.4]
  assign _T_10355 = _T_10353 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31001.4]
  assign _T_10357 = _T_10347 + _T_10352; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31003.4]
  assign _T_10358 = _T_10357 - _T_10355; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31004.4]
  assign _T_10359 = $unsigned(_T_10358); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31005.4]
  assign _T_10360 = _T_10359[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31006.4]
  assign _T_10361 = _T_10355 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31008.4]
  assign _T_10363 = _T_10361 | _T_10347; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31010.4]
  assign _T_10365 = _T_10363 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31012.4]
  assign _T_10366 = _T_10365 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31013.4]
  assign _T_10367 = _T_10352 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31018.4]
  assign _T_10368 = _T_10347 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31019.4]
  assign _T_10369 = _T_10367 | _T_10368; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31020.4]
  assign _T_10371 = _T_10369 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31022.4]
  assign _T_10372 = _T_10371 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31023.4]
  assign _T_10383 = _T_2660 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31040.4]
  assign _T_10384 = _T_2920 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31041.4]
  assign _T_10386 = _T_10384 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31043.4]
  assign _T_10388 = _T_10378 + _T_10383; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31045.4]
  assign _T_10389 = _T_10388 - _T_10386; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31046.4]
  assign _T_10390 = $unsigned(_T_10389); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31047.4]
  assign _T_10391 = _T_10390[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31048.4]
  assign _T_10392 = _T_10386 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31050.4]
  assign _T_10394 = _T_10392 | _T_10378; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31052.4]
  assign _T_10396 = _T_10394 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31054.4]
  assign _T_10397 = _T_10396 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31055.4]
  assign _T_10398 = _T_10383 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31060.4]
  assign _T_10399 = _T_10378 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31061.4]
  assign _T_10400 = _T_10398 | _T_10399; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31062.4]
  assign _T_10402 = _T_10400 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31064.4]
  assign _T_10403 = _T_10402 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31065.4]
  assign _T_10414 = _T_2661 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31082.4]
  assign _T_10415 = _T_2921 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31083.4]
  assign _T_10417 = _T_10415 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31085.4]
  assign _T_10419 = _T_10409 + _T_10414; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31087.4]
  assign _T_10420 = _T_10419 - _T_10417; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31088.4]
  assign _T_10421 = $unsigned(_T_10420); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31089.4]
  assign _T_10422 = _T_10421[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31090.4]
  assign _T_10423 = _T_10417 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31092.4]
  assign _T_10425 = _T_10423 | _T_10409; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31094.4]
  assign _T_10427 = _T_10425 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31096.4]
  assign _T_10428 = _T_10427 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31097.4]
  assign _T_10429 = _T_10414 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31102.4]
  assign _T_10430 = _T_10409 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31103.4]
  assign _T_10431 = _T_10429 | _T_10430; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31104.4]
  assign _T_10433 = _T_10431 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31106.4]
  assign _T_10434 = _T_10433 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31107.4]
  assign _T_10445 = _T_2662 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31124.4]
  assign _T_10446 = _T_2922 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31125.4]
  assign _T_10448 = _T_10446 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31127.4]
  assign _T_10450 = _T_10440 + _T_10445; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31129.4]
  assign _T_10451 = _T_10450 - _T_10448; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31130.4]
  assign _T_10452 = $unsigned(_T_10451); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31131.4]
  assign _T_10453 = _T_10452[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31132.4]
  assign _T_10454 = _T_10448 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31134.4]
  assign _T_10456 = _T_10454 | _T_10440; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31136.4]
  assign _T_10458 = _T_10456 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31138.4]
  assign _T_10459 = _T_10458 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31139.4]
  assign _T_10460 = _T_10445 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31144.4]
  assign _T_10461 = _T_10440 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31145.4]
  assign _T_10462 = _T_10460 | _T_10461; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31146.4]
  assign _T_10464 = _T_10462 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31148.4]
  assign _T_10465 = _T_10464 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31149.4]
  assign _T_10476 = _T_2663 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31166.4]
  assign _T_10477 = _T_2923 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31167.4]
  assign _T_10479 = _T_10477 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31169.4]
  assign _T_10481 = _T_10471 + _T_10476; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31171.4]
  assign _T_10482 = _T_10481 - _T_10479; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31172.4]
  assign _T_10483 = $unsigned(_T_10482); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31173.4]
  assign _T_10484 = _T_10483[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31174.4]
  assign _T_10485 = _T_10479 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31176.4]
  assign _T_10487 = _T_10485 | _T_10471; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31178.4]
  assign _T_10489 = _T_10487 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31180.4]
  assign _T_10490 = _T_10489 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31181.4]
  assign _T_10491 = _T_10476 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31186.4]
  assign _T_10492 = _T_10471 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31187.4]
  assign _T_10493 = _T_10491 | _T_10492; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31188.4]
  assign _T_10495 = _T_10493 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31190.4]
  assign _T_10496 = _T_10495 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31191.4]
  assign _T_10507 = _T_2664 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31208.4]
  assign _T_10508 = _T_2924 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31209.4]
  assign _T_10510 = _T_10508 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31211.4]
  assign _T_10512 = _T_10502 + _T_10507; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31213.4]
  assign _T_10513 = _T_10512 - _T_10510; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31214.4]
  assign _T_10514 = $unsigned(_T_10513); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31215.4]
  assign _T_10515 = _T_10514[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31216.4]
  assign _T_10516 = _T_10510 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31218.4]
  assign _T_10518 = _T_10516 | _T_10502; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31220.4]
  assign _T_10520 = _T_10518 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31222.4]
  assign _T_10521 = _T_10520 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31223.4]
  assign _T_10522 = _T_10507 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31228.4]
  assign _T_10523 = _T_10502 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31229.4]
  assign _T_10524 = _T_10522 | _T_10523; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31230.4]
  assign _T_10526 = _T_10524 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31232.4]
  assign _T_10527 = _T_10526 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31233.4]
  assign _T_10538 = _T_2665 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31250.4]
  assign _T_10539 = _T_2925 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31251.4]
  assign _T_10541 = _T_10539 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31253.4]
  assign _T_10543 = _T_10533 + _T_10538; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31255.4]
  assign _T_10544 = _T_10543 - _T_10541; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31256.4]
  assign _T_10545 = $unsigned(_T_10544); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31257.4]
  assign _T_10546 = _T_10545[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31258.4]
  assign _T_10547 = _T_10541 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31260.4]
  assign _T_10549 = _T_10547 | _T_10533; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31262.4]
  assign _T_10551 = _T_10549 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31264.4]
  assign _T_10552 = _T_10551 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31265.4]
  assign _T_10553 = _T_10538 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31270.4]
  assign _T_10554 = _T_10533 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31271.4]
  assign _T_10555 = _T_10553 | _T_10554; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31272.4]
  assign _T_10557 = _T_10555 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31274.4]
  assign _T_10558 = _T_10557 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31275.4]
  assign _T_10569 = _T_2666 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31292.4]
  assign _T_10570 = _T_2926 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31293.4]
  assign _T_10572 = _T_10570 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31295.4]
  assign _T_10574 = _T_10564 + _T_10569; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31297.4]
  assign _T_10575 = _T_10574 - _T_10572; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31298.4]
  assign _T_10576 = $unsigned(_T_10575); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31299.4]
  assign _T_10577 = _T_10576[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31300.4]
  assign _T_10578 = _T_10572 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31302.4]
  assign _T_10580 = _T_10578 | _T_10564; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31304.4]
  assign _T_10582 = _T_10580 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31306.4]
  assign _T_10583 = _T_10582 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31307.4]
  assign _T_10584 = _T_10569 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31312.4]
  assign _T_10585 = _T_10564 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31313.4]
  assign _T_10586 = _T_10584 | _T_10585; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31314.4]
  assign _T_10588 = _T_10586 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31316.4]
  assign _T_10589 = _T_10588 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31317.4]
  assign _T_10600 = _T_2667 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31334.4]
  assign _T_10601 = _T_2927 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31335.4]
  assign _T_10603 = _T_10601 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31337.4]
  assign _T_10605 = _T_10595 + _T_10600; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31339.4]
  assign _T_10606 = _T_10605 - _T_10603; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31340.4]
  assign _T_10607 = $unsigned(_T_10606); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31341.4]
  assign _T_10608 = _T_10607[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31342.4]
  assign _T_10609 = _T_10603 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31344.4]
  assign _T_10611 = _T_10609 | _T_10595; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31346.4]
  assign _T_10613 = _T_10611 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31348.4]
  assign _T_10614 = _T_10613 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31349.4]
  assign _T_10615 = _T_10600 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31354.4]
  assign _T_10616 = _T_10595 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31355.4]
  assign _T_10617 = _T_10615 | _T_10616; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31356.4]
  assign _T_10619 = _T_10617 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31358.4]
  assign _T_10620 = _T_10619 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31359.4]
  assign _T_10631 = _T_2668 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31376.4]
  assign _T_10632 = _T_2928 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31377.4]
  assign _T_10634 = _T_10632 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31379.4]
  assign _T_10636 = _T_10626 + _T_10631; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31381.4]
  assign _T_10637 = _T_10636 - _T_10634; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31382.4]
  assign _T_10638 = $unsigned(_T_10637); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31383.4]
  assign _T_10639 = _T_10638[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31384.4]
  assign _T_10640 = _T_10634 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31386.4]
  assign _T_10642 = _T_10640 | _T_10626; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31388.4]
  assign _T_10644 = _T_10642 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31390.4]
  assign _T_10645 = _T_10644 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31391.4]
  assign _T_10646 = _T_10631 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31396.4]
  assign _T_10647 = _T_10626 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31397.4]
  assign _T_10648 = _T_10646 | _T_10647; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31398.4]
  assign _T_10650 = _T_10648 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31400.4]
  assign _T_10651 = _T_10650 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31401.4]
  assign _T_10662 = _T_2669 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31418.4]
  assign _T_10663 = _T_2929 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31419.4]
  assign _T_10665 = _T_10663 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31421.4]
  assign _T_10667 = _T_10657 + _T_10662; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31423.4]
  assign _T_10668 = _T_10667 - _T_10665; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31424.4]
  assign _T_10669 = $unsigned(_T_10668); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31425.4]
  assign _T_10670 = _T_10669[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31426.4]
  assign _T_10671 = _T_10665 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31428.4]
  assign _T_10673 = _T_10671 | _T_10657; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31430.4]
  assign _T_10675 = _T_10673 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31432.4]
  assign _T_10676 = _T_10675 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31433.4]
  assign _T_10677 = _T_10662 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31438.4]
  assign _T_10678 = _T_10657 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31439.4]
  assign _T_10679 = _T_10677 | _T_10678; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31440.4]
  assign _T_10681 = _T_10679 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31442.4]
  assign _T_10682 = _T_10681 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31443.4]
  assign _T_10693 = _T_2670 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31460.4]
  assign _T_10694 = _T_2930 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31461.4]
  assign _T_10696 = _T_10694 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31463.4]
  assign _T_10698 = _T_10688 + _T_10693; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31465.4]
  assign _T_10699 = _T_10698 - _T_10696; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31466.4]
  assign _T_10700 = $unsigned(_T_10699); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31467.4]
  assign _T_10701 = _T_10700[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31468.4]
  assign _T_10702 = _T_10696 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31470.4]
  assign _T_10704 = _T_10702 | _T_10688; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31472.4]
  assign _T_10706 = _T_10704 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31474.4]
  assign _T_10707 = _T_10706 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31475.4]
  assign _T_10708 = _T_10693 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31480.4]
  assign _T_10709 = _T_10688 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31481.4]
  assign _T_10710 = _T_10708 | _T_10709; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31482.4]
  assign _T_10712 = _T_10710 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31484.4]
  assign _T_10713 = _T_10712 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31485.4]
  assign _T_10724 = _T_2671 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31502.4]
  assign _T_10725 = _T_2931 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31503.4]
  assign _T_10727 = _T_10725 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31505.4]
  assign _T_10729 = _T_10719 + _T_10724; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31507.4]
  assign _T_10730 = _T_10729 - _T_10727; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31508.4]
  assign _T_10731 = $unsigned(_T_10730); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31509.4]
  assign _T_10732 = _T_10731[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31510.4]
  assign _T_10733 = _T_10727 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31512.4]
  assign _T_10735 = _T_10733 | _T_10719; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31514.4]
  assign _T_10737 = _T_10735 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31516.4]
  assign _T_10738 = _T_10737 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31517.4]
  assign _T_10739 = _T_10724 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31522.4]
  assign _T_10740 = _T_10719 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31523.4]
  assign _T_10741 = _T_10739 | _T_10740; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31524.4]
  assign _T_10743 = _T_10741 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31526.4]
  assign _T_10744 = _T_10743 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31527.4]
  assign _T_10755 = _T_2672 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31544.4]
  assign _T_10756 = _T_2932 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31545.4]
  assign _T_10758 = _T_10756 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31547.4]
  assign _T_10760 = _T_10750 + _T_10755; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31549.4]
  assign _T_10761 = _T_10760 - _T_10758; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31550.4]
  assign _T_10762 = $unsigned(_T_10761); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31551.4]
  assign _T_10763 = _T_10762[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31552.4]
  assign _T_10764 = _T_10758 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31554.4]
  assign _T_10766 = _T_10764 | _T_10750; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31556.4]
  assign _T_10768 = _T_10766 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31558.4]
  assign _T_10769 = _T_10768 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31559.4]
  assign _T_10770 = _T_10755 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31564.4]
  assign _T_10771 = _T_10750 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31565.4]
  assign _T_10772 = _T_10770 | _T_10771; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31566.4]
  assign _T_10774 = _T_10772 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31568.4]
  assign _T_10775 = _T_10774 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31569.4]
  assign _T_10786 = _T_2673 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31586.4]
  assign _T_10787 = _T_2933 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31587.4]
  assign _T_10789 = _T_10787 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31589.4]
  assign _T_10791 = _T_10781 + _T_10786; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31591.4]
  assign _T_10792 = _T_10791 - _T_10789; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31592.4]
  assign _T_10793 = $unsigned(_T_10792); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31593.4]
  assign _T_10794 = _T_10793[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31594.4]
  assign _T_10795 = _T_10789 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31596.4]
  assign _T_10797 = _T_10795 | _T_10781; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31598.4]
  assign _T_10799 = _T_10797 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31600.4]
  assign _T_10800 = _T_10799 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31601.4]
  assign _T_10801 = _T_10786 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31606.4]
  assign _T_10802 = _T_10781 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31607.4]
  assign _T_10803 = _T_10801 | _T_10802; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31608.4]
  assign _T_10805 = _T_10803 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31610.4]
  assign _T_10806 = _T_10805 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31611.4]
  assign _T_10817 = _T_2674 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31628.4]
  assign _T_10818 = _T_2934 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31629.4]
  assign _T_10820 = _T_10818 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31631.4]
  assign _T_10822 = _T_10812 + _T_10817; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31633.4]
  assign _T_10823 = _T_10822 - _T_10820; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31634.4]
  assign _T_10824 = $unsigned(_T_10823); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31635.4]
  assign _T_10825 = _T_10824[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31636.4]
  assign _T_10826 = _T_10820 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31638.4]
  assign _T_10828 = _T_10826 | _T_10812; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31640.4]
  assign _T_10830 = _T_10828 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31642.4]
  assign _T_10831 = _T_10830 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31643.4]
  assign _T_10832 = _T_10817 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31648.4]
  assign _T_10833 = _T_10812 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31649.4]
  assign _T_10834 = _T_10832 | _T_10833; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31650.4]
  assign _T_10836 = _T_10834 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31652.4]
  assign _T_10837 = _T_10836 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31653.4]
  assign _T_10848 = _T_2675 & _T_2942; // @[ToAXI4.scala 229:22:boom.system.TestHarness.MegaBoomConfig.fir@31670.4]
  assign _T_10849 = _T_2935 & _T_2936; // @[ToAXI4.scala 230:22:boom.system.TestHarness.MegaBoomConfig.fir@31671.4]
  assign _T_10851 = _T_10849 & _T_2945; // @[ToAXI4.scala 230:32:boom.system.TestHarness.MegaBoomConfig.fir@31673.4]
  assign _T_10853 = _T_10843 + _T_10848; // @[ToAXI4.scala 231:24:boom.system.TestHarness.MegaBoomConfig.fir@31675.4]
  assign _T_10854 = _T_10853 - _T_10851; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31676.4]
  assign _T_10855 = $unsigned(_T_10854); // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31677.4]
  assign _T_10856 = _T_10855[0:0]; // @[ToAXI4.scala 231:37:boom.system.TestHarness.MegaBoomConfig.fir@31678.4]
  assign _T_10857 = _T_10851 == 1'h0; // @[ToAXI4.scala 233:17:boom.system.TestHarness.MegaBoomConfig.fir@31680.4]
  assign _T_10859 = _T_10857 | _T_10843; // @[ToAXI4.scala 233:22:boom.system.TestHarness.MegaBoomConfig.fir@31682.4]
  assign _T_10861 = _T_10859 | reset; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31684.4]
  assign _T_10862 = _T_10861 == 1'h0; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31685.4]
  assign _T_10863 = _T_10848 == 1'h0; // @[ToAXI4.scala 234:17:boom.system.TestHarness.MegaBoomConfig.fir@31690.4]
  assign _T_10864 = _T_10843 != 1'h1; // @[ToAXI4.scala 234:31:boom.system.TestHarness.MegaBoomConfig.fir@31691.4]
  assign _T_10865 = _T_10863 | _T_10864; // @[ToAXI4.scala 234:22:boom.system.TestHarness.MegaBoomConfig.fir@31692.4]
  assign _T_10867 = _T_10865 | reset; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31694.4]
  assign _T_10868 = _T_10867 == 1'h0; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31695.4]
  assign auto_in_a_ready = _T_2378 & _T_2381; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19454.4]
  assign auto_in_d_valid = _T_2398 ? auto_out_r_valid : auto_out_b_valid; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19454.4]
  assign auto_in_d_bits_opcode = _T_2398 ? 3'h1 : 3'h0; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19454.4]
  assign auto_in_d_bits_size = _T_2398 ? _T_2331 : _T_2333; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19454.4]
  assign auto_in_d_bits_source = _T_2398 ? _T_2330 : _T_2332; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19454.4]
  assign auto_in_d_bits_denied = _T_2398 ? _GEN_516 : _T_2410; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19454.4]
  assign auto_in_d_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19454.4]
  assign auto_in_d_bits_corrupt = _T_2398 ? _T_2411 : 1'h0; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@19454.4]
  assign auto_out_aw_valid = _T_2356_valid & _T_2356_bits_wen; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_id = Queue_1_io_deq_bits_id; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_addr = Queue_1_io_deq_bits_addr; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_len = Queue_1_io_deq_bits_len; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_size = Queue_1_io_deq_bits_size; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_burst = Queue_1_io_deq_bits_burst; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_lock = Queue_1_io_deq_bits_lock; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_cache = Queue_1_io_deq_bits_cache; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_prot = Queue_1_io_deq_bits_prot; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_qos = Queue_1_io_deq_bits_qos; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_aw_bits_user = Queue_1_io_deq_bits_user; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_w_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_w_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_w_bits_strb = Queue_io_deq_bits_strb; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_w_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_b_ready = auto_in_d_ready & _T_2399; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_valid = _T_2356_valid & _T_2360; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_id = Queue_1_io_deq_bits_id; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_addr = Queue_1_io_deq_bits_addr; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_len = Queue_1_io_deq_bits_len; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_size = Queue_1_io_deq_bits_size; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_burst = Queue_1_io_deq_bits_burst; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_lock = Queue_1_io_deq_bits_lock; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_cache = Queue_1_io_deq_bits_cache; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_prot = Queue_1_io_deq_bits_prot; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_qos = Queue_1_io_deq_bits_qos; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_ar_bits_user = Queue_1_io_deq_bits_user; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign auto_out_r_ready = auto_in_d_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@19453.4]
  assign Queue_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@20286.4]
  assign Queue_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@20287.4]
  assign Queue_io_enq_valid = _T_2391 & _T_2379; // @[Decoupled.scala 294:22:boom.system.TestHarness.MegaBoomConfig.fir@20288.4]
  assign Queue_io_enq_bits_data = auto_in_a_bits_data; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20291.4]
  assign Queue_io_enq_bits_strb = auto_in_a_bits_mask; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20290.4]
  assign Queue_io_enq_bits_last = _T_2312 | _T_2313; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20289.4]
  assign Queue_io_deq_ready = auto_out_w_ready; // @[Decoupled.scala 317:15:boom.system.TestHarness.MegaBoomConfig.fir@20298.4]
  assign Queue_1_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@20301.4]
  assign Queue_1_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@20302.4]
  assign Queue_1_io_enq_valid = _T_2384 & _T_2387; // @[Decoupled.scala 294:22:boom.system.TestHarness.MegaBoomConfig.fir@20303.4]
  assign Queue_1_io_enq_bits_id = 8'hff == auto_in_a_bits_source ? 8'hff : _GEN_256; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20314.4]
  assign Queue_1_io_enq_bits_addr = auto_in_a_bits_address; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20313.4]
  assign Queue_1_io_enq_bits_len = _T_2372[10:3]; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20312.4]
  assign Queue_1_io_enq_bits_size = _T_2374 ? 3'h3 : auto_in_a_bits_size; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20311.4]
  assign Queue_1_io_enq_bits_user = {{1'd0}, _T_2329}; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20305.4]
  assign Queue_1_io_enq_bits_wen = _T_2295 == 1'h0; // @[Decoupled.scala 295:21:boom.system.TestHarness.MegaBoomConfig.fir@20304.4]
  assign Queue_1_io_deq_ready = _T_2356_bits_wen ? auto_out_aw_ready : auto_out_ar_ready; // @[Decoupled.scala 317:15:boom.system.TestHarness.MegaBoomConfig.fir@20329.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10843 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_10812 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_10781 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_10750 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_10719 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_10688 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_10657 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_10626 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_10595 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_10564 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10533 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_10502 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_10471 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_10440 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_10409 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_10378 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_10347 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_10316 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_10285 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_10254 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_10223 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_10192 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_10161 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_10130 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_10099 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_10068 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_10037 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_10006 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_9975 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_9944 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_9913 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_9882 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_9851 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_9820 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_9789 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_9758 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_9727 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_9696 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_9665 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_9634 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_9603 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_9572 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_9541 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_9510 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_9479 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_9448 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_9417 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_9386 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_9355 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_9324 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_9293 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_9262 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_9231 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_9200 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_9169 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_9138 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_9107 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_9076 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_9045 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_9014 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_8983 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_8952 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_8921 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_8890 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_8859 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_8828 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_8797 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_8766 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_8735 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_8704 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_8673 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_8642 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_8611 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_8580 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_8549 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_8518 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_8487 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_8456 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_8425 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_8394 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_8363 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_8332 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_8301 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_8270 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_8239 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_8208 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_8177 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_8146 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_8115 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_8084 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_8053 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_8022 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_7991 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_7960 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_7929 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_7898 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_7867 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_7836 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_7805 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_7774 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_7743 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_7712 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_7681 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_7650 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_7619 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_7588 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_7557 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_7526 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_7495 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_7464 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_7433 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_7402 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_7371 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_7340 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_7309 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_7278 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_7247 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_7216 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_7185 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_7154 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_7123 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_7092 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_7061 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_7030 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_6999 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_6968 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_6937 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_6906 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_6875 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_6844 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_6813 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_6782 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_6751 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_6720 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_6689 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_6658 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_6627 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_6596 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_6565 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_6534 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_6503 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_6472 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_6441 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_6410 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_6379 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_6348 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_6317 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_6286 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_6255 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_6224 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_6193 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_6162 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_6131 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_6100 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_6069 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_6038 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_6007 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_5976 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_5945 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_5914 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_5883 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_5852 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_5821 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_5790 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_5759 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_5728 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_5697 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_5666 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_5635 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_5604 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_5573 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_5542 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_5511 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_5480 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_5449 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_5418 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_5387 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_5356 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_5325 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_5294 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_5263 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_5232 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_5201 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_5170 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_5139 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_5108 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_5077 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_5046 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_5015 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_4984 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_4953 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_4922 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_4891 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_4860 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_4829 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_4798 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_4767 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_4736 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_4705 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_4674 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_4643 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_4612 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_4581 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_4550 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_4519 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_4488 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_4457 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_4426 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_4395 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_4364 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_4333 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_4302 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_4271 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_4240 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_4209 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_4178 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_4147 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_4116 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_4085 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_4054 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_4023 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_3992 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_3961 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_3930 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_3899 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_3868 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_3837 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_3806 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_3775 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_3744 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_3713 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_3682 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_3651 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_3620 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_3589 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_3558 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_3527 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_3496 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_3465 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3434 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3403 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3372 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3341 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3310 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3279 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3248 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3217 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3186 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3155 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3124 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3093 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3062 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3031 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3000 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_2969 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_2938 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_2307 = _RAND_256[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_2365 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_2395 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_2403 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_2407 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_10843 <= 1'h0;
    end else begin
      _T_10843 <= _T_10856;
    end
    if (reset) begin
      _T_10812 <= 1'h0;
    end else begin
      _T_10812 <= _T_10825;
    end
    if (reset) begin
      _T_10781 <= 1'h0;
    end else begin
      _T_10781 <= _T_10794;
    end
    if (reset) begin
      _T_10750 <= 1'h0;
    end else begin
      _T_10750 <= _T_10763;
    end
    if (reset) begin
      _T_10719 <= 1'h0;
    end else begin
      _T_10719 <= _T_10732;
    end
    if (reset) begin
      _T_10688 <= 1'h0;
    end else begin
      _T_10688 <= _T_10701;
    end
    if (reset) begin
      _T_10657 <= 1'h0;
    end else begin
      _T_10657 <= _T_10670;
    end
    if (reset) begin
      _T_10626 <= 1'h0;
    end else begin
      _T_10626 <= _T_10639;
    end
    if (reset) begin
      _T_10595 <= 1'h0;
    end else begin
      _T_10595 <= _T_10608;
    end
    if (reset) begin
      _T_10564 <= 1'h0;
    end else begin
      _T_10564 <= _T_10577;
    end
    if (reset) begin
      _T_10533 <= 1'h0;
    end else begin
      _T_10533 <= _T_10546;
    end
    if (reset) begin
      _T_10502 <= 1'h0;
    end else begin
      _T_10502 <= _T_10515;
    end
    if (reset) begin
      _T_10471 <= 1'h0;
    end else begin
      _T_10471 <= _T_10484;
    end
    if (reset) begin
      _T_10440 <= 1'h0;
    end else begin
      _T_10440 <= _T_10453;
    end
    if (reset) begin
      _T_10409 <= 1'h0;
    end else begin
      _T_10409 <= _T_10422;
    end
    if (reset) begin
      _T_10378 <= 1'h0;
    end else begin
      _T_10378 <= _T_10391;
    end
    if (reset) begin
      _T_10347 <= 1'h0;
    end else begin
      _T_10347 <= _T_10360;
    end
    if (reset) begin
      _T_10316 <= 1'h0;
    end else begin
      _T_10316 <= _T_10329;
    end
    if (reset) begin
      _T_10285 <= 1'h0;
    end else begin
      _T_10285 <= _T_10298;
    end
    if (reset) begin
      _T_10254 <= 1'h0;
    end else begin
      _T_10254 <= _T_10267;
    end
    if (reset) begin
      _T_10223 <= 1'h0;
    end else begin
      _T_10223 <= _T_10236;
    end
    if (reset) begin
      _T_10192 <= 1'h0;
    end else begin
      _T_10192 <= _T_10205;
    end
    if (reset) begin
      _T_10161 <= 1'h0;
    end else begin
      _T_10161 <= _T_10174;
    end
    if (reset) begin
      _T_10130 <= 1'h0;
    end else begin
      _T_10130 <= _T_10143;
    end
    if (reset) begin
      _T_10099 <= 1'h0;
    end else begin
      _T_10099 <= _T_10112;
    end
    if (reset) begin
      _T_10068 <= 1'h0;
    end else begin
      _T_10068 <= _T_10081;
    end
    if (reset) begin
      _T_10037 <= 1'h0;
    end else begin
      _T_10037 <= _T_10050;
    end
    if (reset) begin
      _T_10006 <= 1'h0;
    end else begin
      _T_10006 <= _T_10019;
    end
    if (reset) begin
      _T_9975 <= 1'h0;
    end else begin
      _T_9975 <= _T_9988;
    end
    if (reset) begin
      _T_9944 <= 1'h0;
    end else begin
      _T_9944 <= _T_9957;
    end
    if (reset) begin
      _T_9913 <= 1'h0;
    end else begin
      _T_9913 <= _T_9926;
    end
    if (reset) begin
      _T_9882 <= 1'h0;
    end else begin
      _T_9882 <= _T_9895;
    end
    if (reset) begin
      _T_9851 <= 1'h0;
    end else begin
      _T_9851 <= _T_9864;
    end
    if (reset) begin
      _T_9820 <= 1'h0;
    end else begin
      _T_9820 <= _T_9833;
    end
    if (reset) begin
      _T_9789 <= 1'h0;
    end else begin
      _T_9789 <= _T_9802;
    end
    if (reset) begin
      _T_9758 <= 1'h0;
    end else begin
      _T_9758 <= _T_9771;
    end
    if (reset) begin
      _T_9727 <= 1'h0;
    end else begin
      _T_9727 <= _T_9740;
    end
    if (reset) begin
      _T_9696 <= 1'h0;
    end else begin
      _T_9696 <= _T_9709;
    end
    if (reset) begin
      _T_9665 <= 1'h0;
    end else begin
      _T_9665 <= _T_9678;
    end
    if (reset) begin
      _T_9634 <= 1'h0;
    end else begin
      _T_9634 <= _T_9647;
    end
    if (reset) begin
      _T_9603 <= 1'h0;
    end else begin
      _T_9603 <= _T_9616;
    end
    if (reset) begin
      _T_9572 <= 1'h0;
    end else begin
      _T_9572 <= _T_9585;
    end
    if (reset) begin
      _T_9541 <= 1'h0;
    end else begin
      _T_9541 <= _T_9554;
    end
    if (reset) begin
      _T_9510 <= 1'h0;
    end else begin
      _T_9510 <= _T_9523;
    end
    if (reset) begin
      _T_9479 <= 1'h0;
    end else begin
      _T_9479 <= _T_9492;
    end
    if (reset) begin
      _T_9448 <= 1'h0;
    end else begin
      _T_9448 <= _T_9461;
    end
    if (reset) begin
      _T_9417 <= 1'h0;
    end else begin
      _T_9417 <= _T_9430;
    end
    if (reset) begin
      _T_9386 <= 1'h0;
    end else begin
      _T_9386 <= _T_9399;
    end
    if (reset) begin
      _T_9355 <= 1'h0;
    end else begin
      _T_9355 <= _T_9368;
    end
    if (reset) begin
      _T_9324 <= 1'h0;
    end else begin
      _T_9324 <= _T_9337;
    end
    if (reset) begin
      _T_9293 <= 1'h0;
    end else begin
      _T_9293 <= _T_9306;
    end
    if (reset) begin
      _T_9262 <= 1'h0;
    end else begin
      _T_9262 <= _T_9275;
    end
    if (reset) begin
      _T_9231 <= 1'h0;
    end else begin
      _T_9231 <= _T_9244;
    end
    if (reset) begin
      _T_9200 <= 1'h0;
    end else begin
      _T_9200 <= _T_9213;
    end
    if (reset) begin
      _T_9169 <= 1'h0;
    end else begin
      _T_9169 <= _T_9182;
    end
    if (reset) begin
      _T_9138 <= 1'h0;
    end else begin
      _T_9138 <= _T_9151;
    end
    if (reset) begin
      _T_9107 <= 1'h0;
    end else begin
      _T_9107 <= _T_9120;
    end
    if (reset) begin
      _T_9076 <= 1'h0;
    end else begin
      _T_9076 <= _T_9089;
    end
    if (reset) begin
      _T_9045 <= 1'h0;
    end else begin
      _T_9045 <= _T_9058;
    end
    if (reset) begin
      _T_9014 <= 1'h0;
    end else begin
      _T_9014 <= _T_9027;
    end
    if (reset) begin
      _T_8983 <= 1'h0;
    end else begin
      _T_8983 <= _T_8996;
    end
    if (reset) begin
      _T_8952 <= 1'h0;
    end else begin
      _T_8952 <= _T_8965;
    end
    if (reset) begin
      _T_8921 <= 1'h0;
    end else begin
      _T_8921 <= _T_8934;
    end
    if (reset) begin
      _T_8890 <= 1'h0;
    end else begin
      _T_8890 <= _T_8903;
    end
    if (reset) begin
      _T_8859 <= 1'h0;
    end else begin
      _T_8859 <= _T_8872;
    end
    if (reset) begin
      _T_8828 <= 1'h0;
    end else begin
      _T_8828 <= _T_8841;
    end
    if (reset) begin
      _T_8797 <= 1'h0;
    end else begin
      _T_8797 <= _T_8810;
    end
    if (reset) begin
      _T_8766 <= 1'h0;
    end else begin
      _T_8766 <= _T_8779;
    end
    if (reset) begin
      _T_8735 <= 1'h0;
    end else begin
      _T_8735 <= _T_8748;
    end
    if (reset) begin
      _T_8704 <= 1'h0;
    end else begin
      _T_8704 <= _T_8717;
    end
    if (reset) begin
      _T_8673 <= 1'h0;
    end else begin
      _T_8673 <= _T_8686;
    end
    if (reset) begin
      _T_8642 <= 1'h0;
    end else begin
      _T_8642 <= _T_8655;
    end
    if (reset) begin
      _T_8611 <= 1'h0;
    end else begin
      _T_8611 <= _T_8624;
    end
    if (reset) begin
      _T_8580 <= 1'h0;
    end else begin
      _T_8580 <= _T_8593;
    end
    if (reset) begin
      _T_8549 <= 1'h0;
    end else begin
      _T_8549 <= _T_8562;
    end
    if (reset) begin
      _T_8518 <= 1'h0;
    end else begin
      _T_8518 <= _T_8531;
    end
    if (reset) begin
      _T_8487 <= 1'h0;
    end else begin
      _T_8487 <= _T_8500;
    end
    if (reset) begin
      _T_8456 <= 1'h0;
    end else begin
      _T_8456 <= _T_8469;
    end
    if (reset) begin
      _T_8425 <= 1'h0;
    end else begin
      _T_8425 <= _T_8438;
    end
    if (reset) begin
      _T_8394 <= 1'h0;
    end else begin
      _T_8394 <= _T_8407;
    end
    if (reset) begin
      _T_8363 <= 1'h0;
    end else begin
      _T_8363 <= _T_8376;
    end
    if (reset) begin
      _T_8332 <= 1'h0;
    end else begin
      _T_8332 <= _T_8345;
    end
    if (reset) begin
      _T_8301 <= 1'h0;
    end else begin
      _T_8301 <= _T_8314;
    end
    if (reset) begin
      _T_8270 <= 1'h0;
    end else begin
      _T_8270 <= _T_8283;
    end
    if (reset) begin
      _T_8239 <= 1'h0;
    end else begin
      _T_8239 <= _T_8252;
    end
    if (reset) begin
      _T_8208 <= 1'h0;
    end else begin
      _T_8208 <= _T_8221;
    end
    if (reset) begin
      _T_8177 <= 1'h0;
    end else begin
      _T_8177 <= _T_8190;
    end
    if (reset) begin
      _T_8146 <= 1'h0;
    end else begin
      _T_8146 <= _T_8159;
    end
    if (reset) begin
      _T_8115 <= 1'h0;
    end else begin
      _T_8115 <= _T_8128;
    end
    if (reset) begin
      _T_8084 <= 1'h0;
    end else begin
      _T_8084 <= _T_8097;
    end
    if (reset) begin
      _T_8053 <= 1'h0;
    end else begin
      _T_8053 <= _T_8066;
    end
    if (reset) begin
      _T_8022 <= 1'h0;
    end else begin
      _T_8022 <= _T_8035;
    end
    if (reset) begin
      _T_7991 <= 1'h0;
    end else begin
      _T_7991 <= _T_8004;
    end
    if (reset) begin
      _T_7960 <= 1'h0;
    end else begin
      _T_7960 <= _T_7973;
    end
    if (reset) begin
      _T_7929 <= 1'h0;
    end else begin
      _T_7929 <= _T_7942;
    end
    if (reset) begin
      _T_7898 <= 1'h0;
    end else begin
      _T_7898 <= _T_7911;
    end
    if (reset) begin
      _T_7867 <= 1'h0;
    end else begin
      _T_7867 <= _T_7880;
    end
    if (reset) begin
      _T_7836 <= 1'h0;
    end else begin
      _T_7836 <= _T_7849;
    end
    if (reset) begin
      _T_7805 <= 1'h0;
    end else begin
      _T_7805 <= _T_7818;
    end
    if (reset) begin
      _T_7774 <= 1'h0;
    end else begin
      _T_7774 <= _T_7787;
    end
    if (reset) begin
      _T_7743 <= 1'h0;
    end else begin
      _T_7743 <= _T_7756;
    end
    if (reset) begin
      _T_7712 <= 1'h0;
    end else begin
      _T_7712 <= _T_7725;
    end
    if (reset) begin
      _T_7681 <= 1'h0;
    end else begin
      _T_7681 <= _T_7694;
    end
    if (reset) begin
      _T_7650 <= 1'h0;
    end else begin
      _T_7650 <= _T_7663;
    end
    if (reset) begin
      _T_7619 <= 1'h0;
    end else begin
      _T_7619 <= _T_7632;
    end
    if (reset) begin
      _T_7588 <= 1'h0;
    end else begin
      _T_7588 <= _T_7601;
    end
    if (reset) begin
      _T_7557 <= 1'h0;
    end else begin
      _T_7557 <= _T_7570;
    end
    if (reset) begin
      _T_7526 <= 1'h0;
    end else begin
      _T_7526 <= _T_7539;
    end
    if (reset) begin
      _T_7495 <= 1'h0;
    end else begin
      _T_7495 <= _T_7508;
    end
    if (reset) begin
      _T_7464 <= 1'h0;
    end else begin
      _T_7464 <= _T_7477;
    end
    if (reset) begin
      _T_7433 <= 1'h0;
    end else begin
      _T_7433 <= _T_7446;
    end
    if (reset) begin
      _T_7402 <= 1'h0;
    end else begin
      _T_7402 <= _T_7415;
    end
    if (reset) begin
      _T_7371 <= 1'h0;
    end else begin
      _T_7371 <= _T_7384;
    end
    if (reset) begin
      _T_7340 <= 1'h0;
    end else begin
      _T_7340 <= _T_7353;
    end
    if (reset) begin
      _T_7309 <= 1'h0;
    end else begin
      _T_7309 <= _T_7322;
    end
    if (reset) begin
      _T_7278 <= 1'h0;
    end else begin
      _T_7278 <= _T_7291;
    end
    if (reset) begin
      _T_7247 <= 1'h0;
    end else begin
      _T_7247 <= _T_7260;
    end
    if (reset) begin
      _T_7216 <= 1'h0;
    end else begin
      _T_7216 <= _T_7229;
    end
    if (reset) begin
      _T_7185 <= 1'h0;
    end else begin
      _T_7185 <= _T_7198;
    end
    if (reset) begin
      _T_7154 <= 1'h0;
    end else begin
      _T_7154 <= _T_7167;
    end
    if (reset) begin
      _T_7123 <= 1'h0;
    end else begin
      _T_7123 <= _T_7136;
    end
    if (reset) begin
      _T_7092 <= 1'h0;
    end else begin
      _T_7092 <= _T_7105;
    end
    if (reset) begin
      _T_7061 <= 1'h0;
    end else begin
      _T_7061 <= _T_7074;
    end
    if (reset) begin
      _T_7030 <= 1'h0;
    end else begin
      _T_7030 <= _T_7043;
    end
    if (reset) begin
      _T_6999 <= 1'h0;
    end else begin
      _T_6999 <= _T_7012;
    end
    if (reset) begin
      _T_6968 <= 1'h0;
    end else begin
      _T_6968 <= _T_6981;
    end
    if (reset) begin
      _T_6937 <= 1'h0;
    end else begin
      _T_6937 <= _T_6950;
    end
    if (reset) begin
      _T_6906 <= 1'h0;
    end else begin
      _T_6906 <= _T_6919;
    end
    if (reset) begin
      _T_6875 <= 1'h0;
    end else begin
      _T_6875 <= _T_6888;
    end
    if (reset) begin
      _T_6844 <= 1'h0;
    end else begin
      _T_6844 <= _T_6857;
    end
    if (reset) begin
      _T_6813 <= 1'h0;
    end else begin
      _T_6813 <= _T_6826;
    end
    if (reset) begin
      _T_6782 <= 1'h0;
    end else begin
      _T_6782 <= _T_6795;
    end
    if (reset) begin
      _T_6751 <= 1'h0;
    end else begin
      _T_6751 <= _T_6764;
    end
    if (reset) begin
      _T_6720 <= 1'h0;
    end else begin
      _T_6720 <= _T_6733;
    end
    if (reset) begin
      _T_6689 <= 1'h0;
    end else begin
      _T_6689 <= _T_6702;
    end
    if (reset) begin
      _T_6658 <= 1'h0;
    end else begin
      _T_6658 <= _T_6671;
    end
    if (reset) begin
      _T_6627 <= 1'h0;
    end else begin
      _T_6627 <= _T_6640;
    end
    if (reset) begin
      _T_6596 <= 1'h0;
    end else begin
      _T_6596 <= _T_6609;
    end
    if (reset) begin
      _T_6565 <= 1'h0;
    end else begin
      _T_6565 <= _T_6578;
    end
    if (reset) begin
      _T_6534 <= 1'h0;
    end else begin
      _T_6534 <= _T_6547;
    end
    if (reset) begin
      _T_6503 <= 1'h0;
    end else begin
      _T_6503 <= _T_6516;
    end
    if (reset) begin
      _T_6472 <= 1'h0;
    end else begin
      _T_6472 <= _T_6485;
    end
    if (reset) begin
      _T_6441 <= 1'h0;
    end else begin
      _T_6441 <= _T_6454;
    end
    if (reset) begin
      _T_6410 <= 1'h0;
    end else begin
      _T_6410 <= _T_6423;
    end
    if (reset) begin
      _T_6379 <= 1'h0;
    end else begin
      _T_6379 <= _T_6392;
    end
    if (reset) begin
      _T_6348 <= 1'h0;
    end else begin
      _T_6348 <= _T_6361;
    end
    if (reset) begin
      _T_6317 <= 1'h0;
    end else begin
      _T_6317 <= _T_6330;
    end
    if (reset) begin
      _T_6286 <= 1'h0;
    end else begin
      _T_6286 <= _T_6299;
    end
    if (reset) begin
      _T_6255 <= 1'h0;
    end else begin
      _T_6255 <= _T_6268;
    end
    if (reset) begin
      _T_6224 <= 1'h0;
    end else begin
      _T_6224 <= _T_6237;
    end
    if (reset) begin
      _T_6193 <= 1'h0;
    end else begin
      _T_6193 <= _T_6206;
    end
    if (reset) begin
      _T_6162 <= 1'h0;
    end else begin
      _T_6162 <= _T_6175;
    end
    if (reset) begin
      _T_6131 <= 1'h0;
    end else begin
      _T_6131 <= _T_6144;
    end
    if (reset) begin
      _T_6100 <= 1'h0;
    end else begin
      _T_6100 <= _T_6113;
    end
    if (reset) begin
      _T_6069 <= 1'h0;
    end else begin
      _T_6069 <= _T_6082;
    end
    if (reset) begin
      _T_6038 <= 1'h0;
    end else begin
      _T_6038 <= _T_6051;
    end
    if (reset) begin
      _T_6007 <= 1'h0;
    end else begin
      _T_6007 <= _T_6020;
    end
    if (reset) begin
      _T_5976 <= 1'h0;
    end else begin
      _T_5976 <= _T_5989;
    end
    if (reset) begin
      _T_5945 <= 1'h0;
    end else begin
      _T_5945 <= _T_5958;
    end
    if (reset) begin
      _T_5914 <= 1'h0;
    end else begin
      _T_5914 <= _T_5927;
    end
    if (reset) begin
      _T_5883 <= 1'h0;
    end else begin
      _T_5883 <= _T_5896;
    end
    if (reset) begin
      _T_5852 <= 1'h0;
    end else begin
      _T_5852 <= _T_5865;
    end
    if (reset) begin
      _T_5821 <= 1'h0;
    end else begin
      _T_5821 <= _T_5834;
    end
    if (reset) begin
      _T_5790 <= 1'h0;
    end else begin
      _T_5790 <= _T_5803;
    end
    if (reset) begin
      _T_5759 <= 1'h0;
    end else begin
      _T_5759 <= _T_5772;
    end
    if (reset) begin
      _T_5728 <= 1'h0;
    end else begin
      _T_5728 <= _T_5741;
    end
    if (reset) begin
      _T_5697 <= 1'h0;
    end else begin
      _T_5697 <= _T_5710;
    end
    if (reset) begin
      _T_5666 <= 1'h0;
    end else begin
      _T_5666 <= _T_5679;
    end
    if (reset) begin
      _T_5635 <= 1'h0;
    end else begin
      _T_5635 <= _T_5648;
    end
    if (reset) begin
      _T_5604 <= 1'h0;
    end else begin
      _T_5604 <= _T_5617;
    end
    if (reset) begin
      _T_5573 <= 1'h0;
    end else begin
      _T_5573 <= _T_5586;
    end
    if (reset) begin
      _T_5542 <= 1'h0;
    end else begin
      _T_5542 <= _T_5555;
    end
    if (reset) begin
      _T_5511 <= 1'h0;
    end else begin
      _T_5511 <= _T_5524;
    end
    if (reset) begin
      _T_5480 <= 1'h0;
    end else begin
      _T_5480 <= _T_5493;
    end
    if (reset) begin
      _T_5449 <= 1'h0;
    end else begin
      _T_5449 <= _T_5462;
    end
    if (reset) begin
      _T_5418 <= 1'h0;
    end else begin
      _T_5418 <= _T_5431;
    end
    if (reset) begin
      _T_5387 <= 1'h0;
    end else begin
      _T_5387 <= _T_5400;
    end
    if (reset) begin
      _T_5356 <= 1'h0;
    end else begin
      _T_5356 <= _T_5369;
    end
    if (reset) begin
      _T_5325 <= 1'h0;
    end else begin
      _T_5325 <= _T_5338;
    end
    if (reset) begin
      _T_5294 <= 1'h0;
    end else begin
      _T_5294 <= _T_5307;
    end
    if (reset) begin
      _T_5263 <= 1'h0;
    end else begin
      _T_5263 <= _T_5276;
    end
    if (reset) begin
      _T_5232 <= 1'h0;
    end else begin
      _T_5232 <= _T_5245;
    end
    if (reset) begin
      _T_5201 <= 1'h0;
    end else begin
      _T_5201 <= _T_5214;
    end
    if (reset) begin
      _T_5170 <= 1'h0;
    end else begin
      _T_5170 <= _T_5183;
    end
    if (reset) begin
      _T_5139 <= 1'h0;
    end else begin
      _T_5139 <= _T_5152;
    end
    if (reset) begin
      _T_5108 <= 1'h0;
    end else begin
      _T_5108 <= _T_5121;
    end
    if (reset) begin
      _T_5077 <= 1'h0;
    end else begin
      _T_5077 <= _T_5090;
    end
    if (reset) begin
      _T_5046 <= 1'h0;
    end else begin
      _T_5046 <= _T_5059;
    end
    if (reset) begin
      _T_5015 <= 1'h0;
    end else begin
      _T_5015 <= _T_5028;
    end
    if (reset) begin
      _T_4984 <= 1'h0;
    end else begin
      _T_4984 <= _T_4997;
    end
    if (reset) begin
      _T_4953 <= 1'h0;
    end else begin
      _T_4953 <= _T_4966;
    end
    if (reset) begin
      _T_4922 <= 1'h0;
    end else begin
      _T_4922 <= _T_4935;
    end
    if (reset) begin
      _T_4891 <= 1'h0;
    end else begin
      _T_4891 <= _T_4904;
    end
    if (reset) begin
      _T_4860 <= 1'h0;
    end else begin
      _T_4860 <= _T_4873;
    end
    if (reset) begin
      _T_4829 <= 1'h0;
    end else begin
      _T_4829 <= _T_4842;
    end
    if (reset) begin
      _T_4798 <= 1'h0;
    end else begin
      _T_4798 <= _T_4811;
    end
    if (reset) begin
      _T_4767 <= 1'h0;
    end else begin
      _T_4767 <= _T_4780;
    end
    if (reset) begin
      _T_4736 <= 1'h0;
    end else begin
      _T_4736 <= _T_4749;
    end
    if (reset) begin
      _T_4705 <= 1'h0;
    end else begin
      _T_4705 <= _T_4718;
    end
    if (reset) begin
      _T_4674 <= 1'h0;
    end else begin
      _T_4674 <= _T_4687;
    end
    if (reset) begin
      _T_4643 <= 1'h0;
    end else begin
      _T_4643 <= _T_4656;
    end
    if (reset) begin
      _T_4612 <= 1'h0;
    end else begin
      _T_4612 <= _T_4625;
    end
    if (reset) begin
      _T_4581 <= 1'h0;
    end else begin
      _T_4581 <= _T_4594;
    end
    if (reset) begin
      _T_4550 <= 1'h0;
    end else begin
      _T_4550 <= _T_4563;
    end
    if (reset) begin
      _T_4519 <= 1'h0;
    end else begin
      _T_4519 <= _T_4532;
    end
    if (reset) begin
      _T_4488 <= 1'h0;
    end else begin
      _T_4488 <= _T_4501;
    end
    if (reset) begin
      _T_4457 <= 1'h0;
    end else begin
      _T_4457 <= _T_4470;
    end
    if (reset) begin
      _T_4426 <= 1'h0;
    end else begin
      _T_4426 <= _T_4439;
    end
    if (reset) begin
      _T_4395 <= 1'h0;
    end else begin
      _T_4395 <= _T_4408;
    end
    if (reset) begin
      _T_4364 <= 1'h0;
    end else begin
      _T_4364 <= _T_4377;
    end
    if (reset) begin
      _T_4333 <= 1'h0;
    end else begin
      _T_4333 <= _T_4346;
    end
    if (reset) begin
      _T_4302 <= 1'h0;
    end else begin
      _T_4302 <= _T_4315;
    end
    if (reset) begin
      _T_4271 <= 1'h0;
    end else begin
      _T_4271 <= _T_4284;
    end
    if (reset) begin
      _T_4240 <= 1'h0;
    end else begin
      _T_4240 <= _T_4253;
    end
    if (reset) begin
      _T_4209 <= 1'h0;
    end else begin
      _T_4209 <= _T_4222;
    end
    if (reset) begin
      _T_4178 <= 1'h0;
    end else begin
      _T_4178 <= _T_4191;
    end
    if (reset) begin
      _T_4147 <= 1'h0;
    end else begin
      _T_4147 <= _T_4160;
    end
    if (reset) begin
      _T_4116 <= 1'h0;
    end else begin
      _T_4116 <= _T_4129;
    end
    if (reset) begin
      _T_4085 <= 1'h0;
    end else begin
      _T_4085 <= _T_4098;
    end
    if (reset) begin
      _T_4054 <= 1'h0;
    end else begin
      _T_4054 <= _T_4067;
    end
    if (reset) begin
      _T_4023 <= 1'h0;
    end else begin
      _T_4023 <= _T_4036;
    end
    if (reset) begin
      _T_3992 <= 1'h0;
    end else begin
      _T_3992 <= _T_4005;
    end
    if (reset) begin
      _T_3961 <= 1'h0;
    end else begin
      _T_3961 <= _T_3974;
    end
    if (reset) begin
      _T_3930 <= 1'h0;
    end else begin
      _T_3930 <= _T_3943;
    end
    if (reset) begin
      _T_3899 <= 1'h0;
    end else begin
      _T_3899 <= _T_3912;
    end
    if (reset) begin
      _T_3868 <= 1'h0;
    end else begin
      _T_3868 <= _T_3881;
    end
    if (reset) begin
      _T_3837 <= 1'h0;
    end else begin
      _T_3837 <= _T_3850;
    end
    if (reset) begin
      _T_3806 <= 1'h0;
    end else begin
      _T_3806 <= _T_3819;
    end
    if (reset) begin
      _T_3775 <= 1'h0;
    end else begin
      _T_3775 <= _T_3788;
    end
    if (reset) begin
      _T_3744 <= 1'h0;
    end else begin
      _T_3744 <= _T_3757;
    end
    if (reset) begin
      _T_3713 <= 1'h0;
    end else begin
      _T_3713 <= _T_3726;
    end
    if (reset) begin
      _T_3682 <= 1'h0;
    end else begin
      _T_3682 <= _T_3695;
    end
    if (reset) begin
      _T_3651 <= 1'h0;
    end else begin
      _T_3651 <= _T_3664;
    end
    if (reset) begin
      _T_3620 <= 1'h0;
    end else begin
      _T_3620 <= _T_3633;
    end
    if (reset) begin
      _T_3589 <= 1'h0;
    end else begin
      _T_3589 <= _T_3602;
    end
    if (reset) begin
      _T_3558 <= 1'h0;
    end else begin
      _T_3558 <= _T_3571;
    end
    if (reset) begin
      _T_3527 <= 1'h0;
    end else begin
      _T_3527 <= _T_3540;
    end
    if (reset) begin
      _T_3496 <= 1'h0;
    end else begin
      _T_3496 <= _T_3509;
    end
    if (reset) begin
      _T_3465 <= 1'h0;
    end else begin
      _T_3465 <= _T_3478;
    end
    if (reset) begin
      _T_3434 <= 1'h0;
    end else begin
      _T_3434 <= _T_3447;
    end
    if (reset) begin
      _T_3403 <= 1'h0;
    end else begin
      _T_3403 <= _T_3416;
    end
    if (reset) begin
      _T_3372 <= 1'h0;
    end else begin
      _T_3372 <= _T_3385;
    end
    if (reset) begin
      _T_3341 <= 1'h0;
    end else begin
      _T_3341 <= _T_3354;
    end
    if (reset) begin
      _T_3310 <= 1'h0;
    end else begin
      _T_3310 <= _T_3323;
    end
    if (reset) begin
      _T_3279 <= 1'h0;
    end else begin
      _T_3279 <= _T_3292;
    end
    if (reset) begin
      _T_3248 <= 1'h0;
    end else begin
      _T_3248 <= _T_3261;
    end
    if (reset) begin
      _T_3217 <= 1'h0;
    end else begin
      _T_3217 <= _T_3230;
    end
    if (reset) begin
      _T_3186 <= 1'h0;
    end else begin
      _T_3186 <= _T_3199;
    end
    if (reset) begin
      _T_3155 <= 1'h0;
    end else begin
      _T_3155 <= _T_3168;
    end
    if (reset) begin
      _T_3124 <= 1'h0;
    end else begin
      _T_3124 <= _T_3137;
    end
    if (reset) begin
      _T_3093 <= 1'h0;
    end else begin
      _T_3093 <= _T_3106;
    end
    if (reset) begin
      _T_3062 <= 1'h0;
    end else begin
      _T_3062 <= _T_3075;
    end
    if (reset) begin
      _T_3031 <= 1'h0;
    end else begin
      _T_3031 <= _T_3044;
    end
    if (reset) begin
      _T_3000 <= 1'h0;
    end else begin
      _T_3000 <= _T_3013;
    end
    if (reset) begin
      _T_2969 <= 1'h0;
    end else begin
      _T_2969 <= _T_2982;
    end
    if (reset) begin
      _T_2938 <= 1'h0;
    end else begin
      _T_2938 <= _T_2951;
    end
    if (reset) begin
      _T_2307 <= 3'h0;
    end else begin
      if (_T_2297) begin
        if (_T_2311) begin
          if (_T_2296) begin
            _T_2307 <= _T_2302;
          end else begin
            _T_2307 <= 3'h0;
          end
        end else begin
          _T_2307 <= _T_2310;
        end
      end
    end
    if (reset) begin
      _T_2365 <= 1'h0;
    end else begin
      if (_T_2297) begin
        _T_2365 <= _T_2367;
      end
    end
    if (reset) begin
      _T_2395 <= 1'h0;
    end else begin
      if (_T_2396) begin
        _T_2395 <= _T_2397;
      end
    end
    if (reset) begin
      _T_2403 <= 1'h1;
    end else begin
      if (_T_2396) begin
        _T_2403 <= auto_out_r_bits_last;
      end
    end
    if (_T_2403) begin
      _T_2407 <= _T_2405;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:125 assert (a_source  < UInt(BigInt(1) << sourceBits))\n"); // @[ToAXI4.scala 125:14:boom.system.TestHarness.MegaBoomConfig.fir@20263.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[ToAXI4.scala 125:14:boom.system.TestHarness.MegaBoomConfig.fir@20264.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:126 assert (a_size    < UInt(BigInt(1) << sizeBits))\n"); // @[ToAXI4.scala 126:14:boom.system.TestHarness.MegaBoomConfig.fir@20271.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[ToAXI4.scala 126:14:boom.system.TestHarness.MegaBoomConfig.fir@20272.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2957) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@20977.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2957) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@20978.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2963) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@20987.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2963) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@20988.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2988) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21019.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2988) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21020.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2994) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21029.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2994) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21030.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3019) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21061.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3019) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21062.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3025) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21071.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3025) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21072.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3050) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21103.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3050) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21104.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3056) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21113.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3056) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21114.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3081) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21145.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3081) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21146.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3087) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21155.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3087) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21156.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3112) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21187.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3112) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21188.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3118) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21197.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3118) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21198.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3143) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21229.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3143) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21230.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3149) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21239.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3149) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21240.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3174) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21271.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3174) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21272.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3180) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21281.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3180) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21282.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3205) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21313.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3205) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21314.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3211) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21323.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3211) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21324.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3236) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21355.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3236) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21356.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3242) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21365.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3242) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21366.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3267) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21397.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3267) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21398.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3273) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21407.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3273) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21408.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3298) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21439.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3298) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21440.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3304) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21449.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3304) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21450.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3329) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21481.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3329) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21482.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3335) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21491.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3335) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21492.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3360) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21523.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3360) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21524.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3366) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21533.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3366) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21534.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3391) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21565.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3391) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21566.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3397) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21575.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3397) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21576.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3422) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21607.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3422) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21608.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3428) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21617.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3428) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21618.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3453) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21649.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3453) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21650.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3459) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21659.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3459) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21660.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3484) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21691.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3484) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21692.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3490) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21701.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3490) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21702.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3515) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21733.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3515) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21734.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3521) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21743.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3521) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21744.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3546) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21775.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3546) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21776.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3552) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21785.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3552) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21786.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3577) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21817.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3577) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21818.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3583) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21827.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3583) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21828.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3608) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21859.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3608) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21860.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3614) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21869.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3614) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21870.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3639) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21901.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3639) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21902.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3645) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21911.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3645) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21912.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3670) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21943.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3670) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21944.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3676) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21953.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3676) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21954.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3701) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21985.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3701) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@21986.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3707) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21995.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3707) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@21996.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3732) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22027.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3732) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22028.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3738) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22037.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3738) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22038.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3763) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22069.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3763) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22070.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3769) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22079.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3769) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22080.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3794) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22111.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3794) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22112.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3800) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22121.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3800) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22122.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3825) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22153.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3825) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22154.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3831) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22163.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3831) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22164.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3856) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22195.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3856) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22196.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3862) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22205.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3862) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22206.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3887) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22237.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3887) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22238.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3893) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22247.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3893) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22248.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3918) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22279.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3918) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22280.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3924) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22289.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3924) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22290.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3949) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22321.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3949) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22322.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3955) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22331.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3955) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22332.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3980) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22363.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3980) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22364.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3986) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22373.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3986) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22374.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4011) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22405.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4011) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22406.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4017) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22415.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4017) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22416.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4042) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22447.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4042) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22448.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4048) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22457.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4048) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22458.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4073) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22489.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4073) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22490.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4079) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22499.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4079) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22500.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22531.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4104) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22532.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4110) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22541.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4110) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22542.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4135) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22573.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4135) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22574.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4141) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22583.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4141) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22584.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4166) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22615.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4166) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22616.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4172) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22625.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4172) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22626.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4197) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22657.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4197) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22658.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4203) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22667.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4203) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22668.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4228) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22699.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4228) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22700.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4234) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22709.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4234) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22710.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4259) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22741.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4259) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22742.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4265) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22751.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4265) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22752.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4290) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22783.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4290) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22784.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4296) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22793.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4296) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22794.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4321) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22825.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4321) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22826.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4327) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22835.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4327) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22836.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4352) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22867.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4352) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22868.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4358) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22877.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4358) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22878.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4383) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22909.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4383) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22910.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4389) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22919.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4389) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22920.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4414) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22951.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4414) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22952.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4420) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22961.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4420) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@22962.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4445) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22993.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4445) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@22994.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4451) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23003.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4451) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23004.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4476) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23035.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4476) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23036.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4482) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23045.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4482) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23046.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4507) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23077.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4507) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23078.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4513) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23087.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4513) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23088.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4538) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23119.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4538) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23120.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4544) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23129.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4544) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23130.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4569) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23161.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4569) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23162.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4575) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23171.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4575) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23172.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4600) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23203.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4600) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23204.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4606) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23213.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4606) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23214.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4631) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23245.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4631) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23246.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4637) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23255.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4637) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23256.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4662) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23287.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4662) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23288.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4668) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23297.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4668) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23298.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4693) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23329.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4693) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23330.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4699) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23339.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4699) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23340.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4724) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23371.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4724) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23372.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4730) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23381.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4730) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23382.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4755) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23413.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4755) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23414.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4761) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23423.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4761) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23424.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4786) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23455.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4786) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23456.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4792) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23465.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4792) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23466.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4817) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23497.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4817) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23498.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4823) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23507.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4823) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23508.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4848) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23539.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4848) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23540.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4854) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23549.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4854) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23550.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4879) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23581.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4879) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23582.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4885) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23591.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4885) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23592.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4910) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23623.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4910) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23624.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4916) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23633.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4916) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23634.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4941) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23665.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4941) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23666.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4947) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23675.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4947) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23676.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4972) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23707.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4972) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23708.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4978) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23717.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4978) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23718.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5003) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23749.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5003) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23750.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5009) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23759.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5009) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23760.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5034) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23791.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5034) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23792.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5040) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23801.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5040) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23802.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5065) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23833.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5065) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23834.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5071) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23843.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5071) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23844.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5096) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23875.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5096) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23876.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5102) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23885.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5102) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23886.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5127) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23917.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5127) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23918.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5133) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23927.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5133) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23928.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5158) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23959.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5158) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@23960.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5164) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23969.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5164) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@23970.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5189) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24001.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5189) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24002.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5195) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24011.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5195) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24012.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5220) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24043.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5220) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24044.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5226) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24053.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5226) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24054.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5251) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24085.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5251) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24086.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5257) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24095.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5257) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24096.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5282) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24127.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5282) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24128.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5288) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24137.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5288) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24138.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5313) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24169.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5313) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24170.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5319) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24179.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5319) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24180.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5344) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24211.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5344) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24212.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5350) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24221.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5350) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24222.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5375) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24253.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5375) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24254.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5381) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24263.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5381) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24264.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5406) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24295.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5406) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24296.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5412) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24305.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5412) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24306.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5437) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24337.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5437) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24338.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5443) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24347.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5443) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24348.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5468) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24379.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5468) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24380.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5474) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24389.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5474) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24390.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5499) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24421.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5499) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24422.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5505) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24431.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5505) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24432.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5530) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24463.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5530) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24464.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5536) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24473.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5536) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24474.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5561) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24505.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5561) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24506.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5567) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24515.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5567) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24516.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5592) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24547.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5592) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24548.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5598) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24557.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5598) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24558.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5623) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24589.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5623) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24590.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5629) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24599.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5629) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24600.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5654) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24631.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5654) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24632.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5660) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24641.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5660) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24642.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5685) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24673.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5685) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24674.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5691) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24683.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5691) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24684.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5716) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24715.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5716) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24716.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5722) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24725.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5722) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24726.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5747) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24757.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5747) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24758.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5753) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24767.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5753) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24768.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5778) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24799.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5778) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24800.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5784) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24809.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5784) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24810.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5809) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24841.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5809) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24842.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5815) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24851.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5815) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24852.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5840) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24883.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5840) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24884.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5846) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24893.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5846) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24894.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5871) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24925.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5871) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24926.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5877) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24935.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5877) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24936.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5902) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24967.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5902) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@24968.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5908) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24977.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5908) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@24978.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5933) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25009.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5933) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25010.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5939) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25019.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5939) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25020.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5964) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25051.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5964) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25052.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5970) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25061.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5970) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25062.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5995) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25093.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5995) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25094.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6001) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25103.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6001) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25104.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6026) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25135.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6026) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25136.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6032) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25145.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6032) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25146.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6057) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25177.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6057) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25178.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6063) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25187.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6063) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25188.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6088) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25219.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6088) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25220.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6094) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25229.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6094) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25230.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6119) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25261.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6119) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25262.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6125) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25271.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6125) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25272.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6150) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25303.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6150) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25304.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6156) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25313.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6156) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25314.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6181) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25345.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6181) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25346.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6187) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25355.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6187) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25356.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6212) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25387.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6212) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25388.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6218) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25397.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6218) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25398.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6243) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25429.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6243) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25430.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6249) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25439.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6249) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25440.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6274) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25471.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6274) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25472.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6280) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25481.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6280) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25482.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6305) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25513.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6305) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25514.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6311) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25523.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6311) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25524.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6336) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25555.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6336) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25556.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6342) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25565.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6342) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25566.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6367) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25597.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6367) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25598.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6373) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25607.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6373) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25608.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6398) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25639.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6398) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25640.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6404) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25649.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6404) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25650.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6429) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25681.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6429) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25682.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6435) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25691.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6435) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25692.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6460) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25723.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6460) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25724.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6466) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25733.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6466) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25734.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6491) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25765.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6491) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25766.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6497) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25775.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6497) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25776.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6522) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25807.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6522) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25808.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6528) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25817.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6528) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25818.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6553) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25849.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6553) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25850.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6559) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25859.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6559) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25860.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6584) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25891.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6584) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25892.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6590) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25901.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6590) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25902.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6615) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25933.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6615) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25934.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6621) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25943.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6621) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25944.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6646) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25975.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6646) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@25976.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6652) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25985.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6652) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@25986.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6677) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26017.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6677) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26018.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6683) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26027.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6683) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26028.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6708) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26059.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6708) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26060.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6714) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26069.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6714) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26070.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6739) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26101.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6739) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26102.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6745) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26111.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6745) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26112.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6770) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26143.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6770) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26144.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6776) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26153.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6776) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26154.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6801) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26185.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6801) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26186.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6807) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26195.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6807) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26196.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6832) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26227.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6832) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26228.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6838) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26237.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6838) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26238.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6863) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26269.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6863) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26270.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6869) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26279.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6869) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26280.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6894) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26311.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6894) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26312.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6900) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26321.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6900) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26322.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6925) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26353.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6925) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26354.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6931) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26363.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6931) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26364.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6956) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26395.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6956) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26396.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6962) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26405.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6962) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26406.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6987) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26437.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6987) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26438.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6993) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26447.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6993) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26448.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7018) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26479.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7018) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26480.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7024) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26489.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7024) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26490.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7049) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26521.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7049) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26522.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7055) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26531.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7055) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26532.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7080) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26563.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7080) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26564.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7086) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26573.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7086) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26574.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7111) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26605.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7111) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26606.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7117) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26615.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7117) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26616.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7142) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26647.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7142) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26648.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7148) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26657.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7148) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26658.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7173) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26689.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7173) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26690.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7179) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26699.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7179) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26700.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7204) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26731.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7204) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26732.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7210) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26741.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7210) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26742.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7235) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26773.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7235) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26774.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7241) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26783.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7241) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26784.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7266) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26815.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7266) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26816.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7272) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26825.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7272) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26826.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7297) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26857.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7297) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26858.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7303) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26867.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7303) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26868.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7328) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26899.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7328) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26900.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7334) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26909.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7334) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26910.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7359) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26941.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7359) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26942.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7365) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26951.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7365) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26952.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7390) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26983.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7390) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@26984.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7396) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26993.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7396) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@26994.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7421) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27025.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7421) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27026.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7427) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27035.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7427) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27036.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7452) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27067.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7452) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27068.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7458) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27077.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7458) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27078.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7483) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27109.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7483) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27110.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7489) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27119.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7489) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27120.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7514) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27151.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7514) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27152.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7520) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27161.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7520) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27162.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7545) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27193.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7545) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27194.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7551) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27203.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7551) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27204.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7576) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27235.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7576) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27236.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7582) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27245.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7582) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27246.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7607) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27277.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7607) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27278.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7613) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27287.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7613) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27288.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7638) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27319.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7638) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27320.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7644) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27329.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7644) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27330.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7669) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27361.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7669) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27362.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7675) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27371.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7675) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27372.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7700) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27403.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7700) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27404.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7706) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27413.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7706) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27414.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7731) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27445.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7731) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27446.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7737) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27455.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7737) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27456.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7762) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27487.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7762) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27488.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7768) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27497.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7768) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27498.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7793) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27529.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7793) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27530.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7799) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27539.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7799) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27540.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7824) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27571.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7824) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27572.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7830) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27581.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7830) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27582.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7855) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27613.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7855) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27614.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7861) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27623.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7861) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27624.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7886) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27655.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7886) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27656.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7892) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27665.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7892) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27666.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7917) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27697.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7917) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27698.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7923) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27707.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7923) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27708.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7948) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27739.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7948) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27740.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7954) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27749.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7954) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27750.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7979) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27781.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7979) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27782.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7985) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27791.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7985) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27792.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8010) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27823.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8010) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27824.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8016) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27833.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8016) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27834.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8041) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27865.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8041) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27866.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8047) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27875.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8047) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27876.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8072) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27907.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8072) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27908.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8078) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27917.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8078) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27918.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8103) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27949.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8103) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27950.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8109) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27959.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8109) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@27960.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8134) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27991.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8134) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@27992.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8140) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28001.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8140) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28002.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8165) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28033.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8165) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28034.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8171) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28043.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8171) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28044.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8196) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28075.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8196) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28076.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8202) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28085.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8202) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28086.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8227) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28117.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8227) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28118.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8233) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28127.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8233) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28128.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8258) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28159.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8258) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28160.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8264) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28169.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8264) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28170.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8289) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28201.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8289) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28202.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8295) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28211.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8295) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28212.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8320) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28243.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8320) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28244.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8326) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28253.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8326) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28254.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8351) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28285.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8351) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28286.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8357) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28295.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8357) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28296.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8382) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28327.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8382) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28328.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8388) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28337.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8388) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28338.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8413) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28369.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8413) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28370.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8419) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28379.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8419) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28380.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8444) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28411.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8444) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28412.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8450) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28421.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8450) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28422.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8475) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28453.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8475) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28454.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8481) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28463.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8481) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28464.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8506) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28495.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8506) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28496.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8512) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28505.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8512) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28506.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8537) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28537.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8537) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28538.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8543) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28547.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8543) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28548.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8568) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28579.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8568) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28580.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8574) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28589.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8574) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28590.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8599) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28621.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8599) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28622.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8605) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28631.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8605) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28632.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8630) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28663.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8630) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28664.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8636) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28673.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8636) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28674.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8661) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28705.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8661) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28706.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8667) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28715.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8667) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28716.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8692) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28747.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8692) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28748.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8698) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28757.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8698) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28758.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8723) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28789.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8723) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28790.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8729) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28799.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8729) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28800.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8754) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28831.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8754) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28832.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8760) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28841.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8760) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28842.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8785) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28873.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8785) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28874.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8791) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28883.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8791) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28884.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8816) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28915.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8816) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28916.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8822) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28925.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8822) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28926.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8847) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28957.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8847) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28958.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8853) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28967.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8853) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@28968.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8878) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@28999.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8878) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29000.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8884) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29009.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8884) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29010.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8909) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29041.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8909) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29042.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8915) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29051.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8915) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29052.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8940) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29083.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8940) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29084.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8946) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29093.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8946) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29094.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8971) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29125.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8971) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29126.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8977) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29135.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8977) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29136.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9002) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29167.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9002) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29168.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9008) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29177.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9008) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29178.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9033) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29209.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9033) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29210.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9039) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29219.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9039) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29220.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9064) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29251.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9064) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29252.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9070) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29261.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9070) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29262.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9095) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29293.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9095) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29294.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9101) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29303.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9101) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29304.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9126) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29335.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9126) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29336.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9132) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29345.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9132) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29346.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9157) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29377.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9157) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29378.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9163) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29387.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9163) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29388.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9188) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29419.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9188) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29420.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9194) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29429.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9194) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29430.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9219) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29461.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9219) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29462.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9225) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29471.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9225) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29472.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9250) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29503.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9250) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29504.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9256) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29513.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9256) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29514.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9281) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29545.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9281) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29546.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9287) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29555.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9287) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29556.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9312) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29587.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9312) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29588.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9318) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29597.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9318) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29598.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9343) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29629.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9343) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29630.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9349) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29639.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9349) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29640.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9374) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29671.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9374) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29672.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9380) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29681.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9380) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29682.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9405) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29713.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9405) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29714.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9411) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29723.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9411) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29724.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9436) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29755.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9436) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29756.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9442) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29765.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9442) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29766.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9467) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29797.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9467) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29798.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9473) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29807.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9473) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29808.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9498) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29839.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9498) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29840.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9504) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29849.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9504) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29850.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9529) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29881.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9529) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29882.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9535) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29891.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9535) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29892.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9560) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29923.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9560) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29924.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9566) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29933.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9566) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29934.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9591) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29965.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9591) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@29966.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9597) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29975.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9597) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@29976.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9622) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30007.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9622) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30008.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9628) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30017.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9628) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30018.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9653) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30049.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9653) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30050.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9659) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30059.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9659) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30060.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9684) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30091.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9684) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30092.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9690) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30101.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9690) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30102.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9715) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30133.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9715) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30134.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9721) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30143.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9721) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30144.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9746) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30175.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9746) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30176.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9752) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30185.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9752) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30186.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9777) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30217.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9777) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30218.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9783) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30227.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9783) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30228.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9808) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30259.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9808) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30260.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9814) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30269.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9814) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30270.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9839) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30301.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9839) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30302.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9845) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30311.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9845) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30312.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9870) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30343.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9870) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30344.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9876) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30353.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9876) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30354.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9901) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30385.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9901) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30386.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9907) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30395.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9907) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30396.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9932) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30427.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9932) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30428.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9938) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30437.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9938) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30438.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9963) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30469.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9963) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30470.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9969) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30479.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9969) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30480.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9994) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30511.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9994) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30512.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10000) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30521.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10000) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30522.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10025) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30553.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10025) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30554.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10031) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30563.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10031) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30564.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10056) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30595.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10056) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30596.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10062) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30605.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10062) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30606.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10087) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30637.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10087) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30638.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10093) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30647.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10093) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30648.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10118) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30679.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10118) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30680.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10124) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30689.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10124) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30690.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10149) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30721.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10149) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30722.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10155) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30731.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10155) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30732.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10180) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30763.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10180) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30764.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10186) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30773.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10186) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30774.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10211) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30805.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10211) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30806.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10217) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30815.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10217) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30816.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10242) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30847.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10242) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30848.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10248) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30857.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10248) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30858.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10273) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30889.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10273) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30890.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10279) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30899.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10279) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30900.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10304) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30931.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10304) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30932.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10310) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30941.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10310) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30942.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10335) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30973.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10335) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@30974.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10341) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30983.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10341) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@30984.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10366) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31015.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10366) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31016.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10372) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31025.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10372) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31026.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10397) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31057.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10397) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31058.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10403) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31067.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10403) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31068.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10428) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31099.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10428) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31100.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10434) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31109.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10434) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31110.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10459) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31141.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10459) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31142.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10465) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31151.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10465) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31152.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10490) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31183.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10490) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31184.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10496) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31193.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10496) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31194.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10521) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31225.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10521) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31226.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10527) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31235.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10527) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31236.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10552) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31267.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10552) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31268.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10558) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31277.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10558) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31278.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10583) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31309.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10583) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31310.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10589) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31319.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10589) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31320.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10614) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31351.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10614) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31352.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10620) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31361.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10620) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31362.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10645) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31393.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10645) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31394.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10651) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31403.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10651) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31404.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10676) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31435.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10676) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31436.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10682) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31445.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10682) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31446.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10707) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31477.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10707) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31478.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10713) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31487.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10713) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31488.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10738) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31519.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10738) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31520.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10744) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31529.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10744) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31530.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10769) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31561.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10769) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31562.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10775) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31571.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10775) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31572.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10800) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31603.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10800) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31604.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10806) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31613.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10806) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31614.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10831) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31645.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10831) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31646.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10837) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31655.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10837) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31656.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10862) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31687.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10862) begin
          $fatal; // @[ToAXI4.scala 233:16:boom.system.TestHarness.MegaBoomConfig.fir@31688.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10868) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31697.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10868) begin
          $fatal; // @[ToAXI4.scala 234:16:boom.system.TestHarness.MegaBoomConfig.fir@31698.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SimMemoryBus( // @[:boom.system.TestHarness.MegaBoomConfig.fir@31735.2] //SimpleLazyModule17
  input         clock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31736.4]
  input         reset, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31737.4]
  output        auto_buffer_in_a_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input         auto_buffer_in_a_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [2:0]  auto_buffer_in_a_bits_opcode, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [2:0]  auto_buffer_in_a_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [7:0]  auto_buffer_in_a_bits_source, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [31:0] auto_buffer_in_a_bits_address, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [7:0]  auto_buffer_in_a_bits_mask, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [63:0] auto_buffer_in_a_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input         auto_buffer_in_d_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_buffer_in_d_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [2:0]  auto_buffer_in_d_bits_opcode, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [1:0]  auto_buffer_in_d_bits_param, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [2:0]  auto_buffer_in_d_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [7:0]  auto_buffer_in_d_bits_source, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_buffer_in_d_bits_denied, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [63:0] auto_buffer_in_d_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_buffer_in_d_bits_corrupt, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input         auto_axi4yank_out_aw_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_axi4yank_out_aw_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [3:0]  auto_axi4yank_out_aw_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [31:0] auto_axi4yank_out_aw_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [7:0]  auto_axi4yank_out_aw_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [2:0]  auto_axi4yank_out_aw_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [1:0]  auto_axi4yank_out_aw_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_axi4yank_out_aw_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [3:0]  auto_axi4yank_out_aw_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [2:0]  auto_axi4yank_out_aw_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [3:0]  auto_axi4yank_out_aw_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input         auto_axi4yank_out_w_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_axi4yank_out_w_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [63:0] auto_axi4yank_out_w_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [7:0]  auto_axi4yank_out_w_bits_strb, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_axi4yank_out_w_bits_last, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_axi4yank_out_b_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input         auto_axi4yank_out_b_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [3:0]  auto_axi4yank_out_b_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [1:0]  auto_axi4yank_out_b_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input         auto_axi4yank_out_ar_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_axi4yank_out_ar_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [3:0]  auto_axi4yank_out_ar_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [31:0] auto_axi4yank_out_ar_bits_addr, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [7:0]  auto_axi4yank_out_ar_bits_len, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [2:0]  auto_axi4yank_out_ar_bits_size, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [1:0]  auto_axi4yank_out_ar_bits_burst, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_axi4yank_out_ar_bits_lock, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [3:0]  auto_axi4yank_out_ar_bits_cache, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [2:0]  auto_axi4yank_out_ar_bits_prot, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output [3:0]  auto_axi4yank_out_ar_bits_qos, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  output        auto_axi4yank_out_r_ready, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input         auto_axi4yank_out_r_valid, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [3:0]  auto_axi4yank_out_r_bits_id, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [63:0] auto_axi4yank_out_r_bits_data, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input  [1:0]  auto_axi4yank_out_r_bits_resp, // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
  input         auto_axi4yank_out_r_bits_last // @[:boom.system.TestHarness.MegaBoomConfig.fir@31738.4]
);
  wire  axi4yank_clock; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_reset; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_aw_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_aw_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_in_aw_bits_id; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [31:0] axi4yank_auto_in_aw_bits_addr; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [7:0] axi4yank_auto_in_aw_bits_len; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [2:0] axi4yank_auto_in_aw_bits_size; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [1:0] axi4yank_auto_in_aw_bits_burst; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_aw_bits_lock; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_in_aw_bits_cache; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [2:0] axi4yank_auto_in_aw_bits_prot; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_in_aw_bits_qos; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [15:0] axi4yank_auto_in_aw_bits_user; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_w_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_w_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [63:0] axi4yank_auto_in_w_bits_data; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [7:0] axi4yank_auto_in_w_bits_strb; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_w_bits_last; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_b_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_b_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_in_b_bits_id; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [1:0] axi4yank_auto_in_b_bits_resp; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [15:0] axi4yank_auto_in_b_bits_user; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_ar_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_ar_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_in_ar_bits_id; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [31:0] axi4yank_auto_in_ar_bits_addr; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [7:0] axi4yank_auto_in_ar_bits_len; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [2:0] axi4yank_auto_in_ar_bits_size; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [1:0] axi4yank_auto_in_ar_bits_burst; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_ar_bits_lock; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_in_ar_bits_cache; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [2:0] axi4yank_auto_in_ar_bits_prot; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_in_ar_bits_qos; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [15:0] axi4yank_auto_in_ar_bits_user; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_r_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_r_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_in_r_bits_id; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [63:0] axi4yank_auto_in_r_bits_data; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [1:0] axi4yank_auto_in_r_bits_resp; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [15:0] axi4yank_auto_in_r_bits_user; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_in_r_bits_last; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_aw_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_aw_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_out_aw_bits_id; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [31:0] axi4yank_auto_out_aw_bits_addr; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [7:0] axi4yank_auto_out_aw_bits_len; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [2:0] axi4yank_auto_out_aw_bits_size; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [1:0] axi4yank_auto_out_aw_bits_burst; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_aw_bits_lock; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_out_aw_bits_cache; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [2:0] axi4yank_auto_out_aw_bits_prot; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_out_aw_bits_qos; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_w_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_w_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [63:0] axi4yank_auto_out_w_bits_data; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [7:0] axi4yank_auto_out_w_bits_strb; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_w_bits_last; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_b_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_b_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_out_b_bits_id; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [1:0] axi4yank_auto_out_b_bits_resp; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_ar_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_ar_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_out_ar_bits_id; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [31:0] axi4yank_auto_out_ar_bits_addr; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [7:0] axi4yank_auto_out_ar_bits_len; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [2:0] axi4yank_auto_out_ar_bits_size; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [1:0] axi4yank_auto_out_ar_bits_burst; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_ar_bits_lock; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_out_ar_bits_cache; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [2:0] axi4yank_auto_out_ar_bits_prot; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_out_ar_bits_qos; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_r_ready; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_r_valid; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [3:0] axi4yank_auto_out_r_bits_id; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [63:0] axi4yank_auto_out_r_bits_data; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire [1:0] axi4yank_auto_out_r_bits_resp; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4yank_auto_out_r_bits_last; // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
  wire  axi4index_auto_in_aw_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_aw_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_in_aw_bits_id; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [31:0] axi4index_auto_in_aw_bits_addr; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_in_aw_bits_len; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [2:0] axi4index_auto_in_aw_bits_size; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [1:0] axi4index_auto_in_aw_bits_burst; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_aw_bits_lock; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_in_aw_bits_cache; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [2:0] axi4index_auto_in_aw_bits_prot; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_in_aw_bits_qos; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [11:0] axi4index_auto_in_aw_bits_user; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_w_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_w_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [63:0] axi4index_auto_in_w_bits_data; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_in_w_bits_strb; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_w_bits_last; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_b_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_b_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_in_b_bits_id; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [1:0] axi4index_auto_in_b_bits_resp; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [11:0] axi4index_auto_in_b_bits_user; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_ar_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_ar_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_in_ar_bits_id; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [31:0] axi4index_auto_in_ar_bits_addr; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_in_ar_bits_len; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [2:0] axi4index_auto_in_ar_bits_size; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [1:0] axi4index_auto_in_ar_bits_burst; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_ar_bits_lock; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_in_ar_bits_cache; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [2:0] axi4index_auto_in_ar_bits_prot; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_in_ar_bits_qos; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [11:0] axi4index_auto_in_ar_bits_user; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_r_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_r_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_in_r_bits_id; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [63:0] axi4index_auto_in_r_bits_data; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [1:0] axi4index_auto_in_r_bits_resp; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [11:0] axi4index_auto_in_r_bits_user; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_in_r_bits_last; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_aw_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_aw_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_out_aw_bits_id; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [31:0] axi4index_auto_out_aw_bits_addr; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_out_aw_bits_len; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [2:0] axi4index_auto_out_aw_bits_size; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [1:0] axi4index_auto_out_aw_bits_burst; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_aw_bits_lock; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_out_aw_bits_cache; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [2:0] axi4index_auto_out_aw_bits_prot; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_out_aw_bits_qos; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [15:0] axi4index_auto_out_aw_bits_user; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_w_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_w_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [63:0] axi4index_auto_out_w_bits_data; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_out_w_bits_strb; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_w_bits_last; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_b_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_b_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_out_b_bits_id; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [1:0] axi4index_auto_out_b_bits_resp; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [15:0] axi4index_auto_out_b_bits_user; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_ar_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_ar_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_out_ar_bits_id; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [31:0] axi4index_auto_out_ar_bits_addr; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [7:0] axi4index_auto_out_ar_bits_len; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [2:0] axi4index_auto_out_ar_bits_size; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [1:0] axi4index_auto_out_ar_bits_burst; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_ar_bits_lock; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_out_ar_bits_cache; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [2:0] axi4index_auto_out_ar_bits_prot; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_out_ar_bits_qos; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [15:0] axi4index_auto_out_ar_bits_user; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_r_ready; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_r_valid; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [3:0] axi4index_auto_out_r_bits_id; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [63:0] axi4index_auto_out_r_bits_data; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [1:0] axi4index_auto_out_r_bits_resp; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire [15:0] axi4index_auto_out_r_bits_user; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  axi4index_auto_out_r_bits_last; // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
  wire  tl2axi4_clock; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_reset; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_in_a_ready; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_in_a_valid; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [2:0] tl2axi4_auto_in_a_bits_opcode; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [2:0] tl2axi4_auto_in_a_bits_size; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_in_a_bits_source; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [31:0] tl2axi4_auto_in_a_bits_address; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_in_a_bits_mask; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [63:0] tl2axi4_auto_in_a_bits_data; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_in_d_ready; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_in_d_valid; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [2:0] tl2axi4_auto_in_d_bits_opcode; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [2:0] tl2axi4_auto_in_d_bits_size; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_in_d_bits_source; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_in_d_bits_denied; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [63:0] tl2axi4_auto_in_d_bits_data; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_in_d_bits_corrupt; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_aw_ready; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_aw_valid; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_out_aw_bits_id; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [31:0] tl2axi4_auto_out_aw_bits_addr; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_out_aw_bits_len; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [2:0] tl2axi4_auto_out_aw_bits_size; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [1:0] tl2axi4_auto_out_aw_bits_burst; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_aw_bits_lock; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [3:0] tl2axi4_auto_out_aw_bits_cache; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [2:0] tl2axi4_auto_out_aw_bits_prot; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [3:0] tl2axi4_auto_out_aw_bits_qos; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [11:0] tl2axi4_auto_out_aw_bits_user; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_w_ready; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_w_valid; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [63:0] tl2axi4_auto_out_w_bits_data; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_out_w_bits_strb; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_w_bits_last; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_b_ready; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_b_valid; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_out_b_bits_id; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [1:0] tl2axi4_auto_out_b_bits_resp; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [11:0] tl2axi4_auto_out_b_bits_user; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_ar_ready; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_ar_valid; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_out_ar_bits_id; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [31:0] tl2axi4_auto_out_ar_bits_addr; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_out_ar_bits_len; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [2:0] tl2axi4_auto_out_ar_bits_size; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [1:0] tl2axi4_auto_out_ar_bits_burst; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_ar_bits_lock; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [3:0] tl2axi4_auto_out_ar_bits_cache; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [2:0] tl2axi4_auto_out_ar_bits_prot; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [3:0] tl2axi4_auto_out_ar_bits_qos; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [11:0] tl2axi4_auto_out_ar_bits_user; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_r_ready; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_r_valid; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [7:0] tl2axi4_auto_out_r_bits_id; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [63:0] tl2axi4_auto_out_r_bits_data; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [1:0] tl2axi4_auto_out_r_bits_resp; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire [11:0] tl2axi4_auto_out_r_bits_user; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  tl2axi4_auto_out_r_bits_last; // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [2:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [7:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [31:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [1:0] buffer_auto_in_d_bits_param; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [2:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [7:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [2:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [7:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [31:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [1:0] buffer_auto_out_d_bits_param; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [2:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [7:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_out_d_bits_denied; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  wire  buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
  AXI4UserYanker_2 axi4yank ( // @[UserYanker.scala 96:30:boom.system.TestHarness.MegaBoomConfig.fir@31743.4]
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_aw_ready(axi4yank_auto_in_aw_ready),
    .auto_in_aw_valid(axi4yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4yank_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4yank_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4yank_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4yank_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4yank_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4yank_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(axi4yank_auto_in_aw_bits_user),
    .auto_in_w_ready(axi4yank_auto_in_w_ready),
    .auto_in_w_valid(axi4yank_auto_in_w_valid),
    .auto_in_w_bits_data(axi4yank_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4yank_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4yank_auto_in_w_bits_last),
    .auto_in_b_ready(axi4yank_auto_in_b_ready),
    .auto_in_b_valid(axi4yank_auto_in_b_valid),
    .auto_in_b_bits_id(axi4yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4yank_auto_in_b_bits_resp),
    .auto_in_b_bits_user(axi4yank_auto_in_b_bits_user),
    .auto_in_ar_ready(axi4yank_auto_in_ar_ready),
    .auto_in_ar_valid(axi4yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4yank_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4yank_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4yank_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4yank_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4yank_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4yank_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(axi4yank_auto_in_ar_bits_user),
    .auto_in_r_ready(axi4yank_auto_in_r_ready),
    .auto_in_r_valid(axi4yank_auto_in_r_valid),
    .auto_in_r_bits_id(axi4yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4yank_auto_in_r_bits_resp),
    .auto_in_r_bits_user(axi4yank_auto_in_r_bits_user),
    .auto_in_r_bits_last(axi4yank_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4yank_auto_out_aw_ready),
    .auto_out_aw_valid(axi4yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4yank_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4yank_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4yank_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4yank_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4yank_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4yank_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4yank_auto_out_aw_bits_qos),
    .auto_out_w_ready(axi4yank_auto_out_w_ready),
    .auto_out_w_valid(axi4yank_auto_out_w_valid),
    .auto_out_w_bits_data(axi4yank_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4yank_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4yank_auto_out_w_bits_last),
    .auto_out_b_ready(axi4yank_auto_out_b_ready),
    .auto_out_b_valid(axi4yank_auto_out_b_valid),
    .auto_out_b_bits_id(axi4yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4yank_auto_out_ar_ready),
    .auto_out_ar_valid(axi4yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4yank_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4yank_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4yank_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4yank_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4yank_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4yank_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4yank_auto_out_ar_bits_qos),
    .auto_out_r_ready(axi4yank_auto_out_r_ready),
    .auto_out_r_valid(axi4yank_auto_out_r_valid),
    .auto_out_r_bits_id(axi4yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4yank_auto_out_r_bits_last)
  );
  AXI4IdIndexer_2 axi4index ( // @[IdIndexer.scala 80:31:boom.system.TestHarness.MegaBoomConfig.fir@31749.4]
    .auto_in_aw_ready(axi4index_auto_in_aw_ready),
    .auto_in_aw_valid(axi4index_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4index_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4index_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4index_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4index_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4index_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4index_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4index_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4index_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4index_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(axi4index_auto_in_aw_bits_user),
    .auto_in_w_ready(axi4index_auto_in_w_ready),
    .auto_in_w_valid(axi4index_auto_in_w_valid),
    .auto_in_w_bits_data(axi4index_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4index_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4index_auto_in_w_bits_last),
    .auto_in_b_ready(axi4index_auto_in_b_ready),
    .auto_in_b_valid(axi4index_auto_in_b_valid),
    .auto_in_b_bits_id(axi4index_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4index_auto_in_b_bits_resp),
    .auto_in_b_bits_user(axi4index_auto_in_b_bits_user),
    .auto_in_ar_ready(axi4index_auto_in_ar_ready),
    .auto_in_ar_valid(axi4index_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4index_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4index_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4index_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4index_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4index_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4index_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4index_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4index_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4index_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(axi4index_auto_in_ar_bits_user),
    .auto_in_r_ready(axi4index_auto_in_r_ready),
    .auto_in_r_valid(axi4index_auto_in_r_valid),
    .auto_in_r_bits_id(axi4index_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4index_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4index_auto_in_r_bits_resp),
    .auto_in_r_bits_user(axi4index_auto_in_r_bits_user),
    .auto_in_r_bits_last(axi4index_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4index_auto_out_aw_ready),
    .auto_out_aw_valid(axi4index_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4index_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4index_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4index_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4index_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4index_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4index_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4index_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4index_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4index_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(axi4index_auto_out_aw_bits_user),
    .auto_out_w_ready(axi4index_auto_out_w_ready),
    .auto_out_w_valid(axi4index_auto_out_w_valid),
    .auto_out_w_bits_data(axi4index_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4index_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4index_auto_out_w_bits_last),
    .auto_out_b_ready(axi4index_auto_out_b_ready),
    .auto_out_b_valid(axi4index_auto_out_b_valid),
    .auto_out_b_bits_id(axi4index_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4index_auto_out_b_bits_resp),
    .auto_out_b_bits_user(axi4index_auto_out_b_bits_user),
    .auto_out_ar_ready(axi4index_auto_out_ar_ready),
    .auto_out_ar_valid(axi4index_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4index_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4index_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4index_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4index_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4index_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4index_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4index_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4index_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4index_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(axi4index_auto_out_ar_bits_user),
    .auto_out_r_ready(axi4index_auto_out_r_ready),
    .auto_out_r_valid(axi4index_auto_out_r_valid),
    .auto_out_r_bits_id(axi4index_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4index_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4index_auto_out_r_bits_resp),
    .auto_out_r_bits_user(axi4index_auto_out_r_bits_user),
    .auto_out_r_bits_last(axi4index_auto_out_r_bits_last)
  );
  TLToAXI4_1 tl2axi4 ( // @[ToAXI4.scala 254:29:boom.system.TestHarness.MegaBoomConfig.fir@31755.4]
    .clock(tl2axi4_clock),
    .reset(tl2axi4_reset),
    .auto_in_a_ready(tl2axi4_auto_in_a_ready),
    .auto_in_a_valid(tl2axi4_auto_in_a_valid),
    .auto_in_a_bits_opcode(tl2axi4_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(tl2axi4_auto_in_a_bits_size),
    .auto_in_a_bits_source(tl2axi4_auto_in_a_bits_source),
    .auto_in_a_bits_address(tl2axi4_auto_in_a_bits_address),
    .auto_in_a_bits_mask(tl2axi4_auto_in_a_bits_mask),
    .auto_in_a_bits_data(tl2axi4_auto_in_a_bits_data),
    .auto_in_d_ready(tl2axi4_auto_in_d_ready),
    .auto_in_d_valid(tl2axi4_auto_in_d_valid),
    .auto_in_d_bits_opcode(tl2axi4_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(tl2axi4_auto_in_d_bits_size),
    .auto_in_d_bits_source(tl2axi4_auto_in_d_bits_source),
    .auto_in_d_bits_denied(tl2axi4_auto_in_d_bits_denied),
    .auto_in_d_bits_data(tl2axi4_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(tl2axi4_auto_in_d_bits_corrupt),
    .auto_out_aw_ready(tl2axi4_auto_out_aw_ready),
    .auto_out_aw_valid(tl2axi4_auto_out_aw_valid),
    .auto_out_aw_bits_id(tl2axi4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(tl2axi4_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(tl2axi4_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(tl2axi4_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(tl2axi4_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(tl2axi4_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(tl2axi4_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(tl2axi4_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(tl2axi4_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(tl2axi4_auto_out_aw_bits_user),
    .auto_out_w_ready(tl2axi4_auto_out_w_ready),
    .auto_out_w_valid(tl2axi4_auto_out_w_valid),
    .auto_out_w_bits_data(tl2axi4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(tl2axi4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(tl2axi4_auto_out_w_bits_last),
    .auto_out_b_ready(tl2axi4_auto_out_b_ready),
    .auto_out_b_valid(tl2axi4_auto_out_b_valid),
    .auto_out_b_bits_id(tl2axi4_auto_out_b_bits_id),
    .auto_out_b_bits_resp(tl2axi4_auto_out_b_bits_resp),
    .auto_out_b_bits_user(tl2axi4_auto_out_b_bits_user),
    .auto_out_ar_ready(tl2axi4_auto_out_ar_ready),
    .auto_out_ar_valid(tl2axi4_auto_out_ar_valid),
    .auto_out_ar_bits_id(tl2axi4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(tl2axi4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(tl2axi4_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(tl2axi4_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(tl2axi4_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(tl2axi4_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(tl2axi4_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(tl2axi4_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(tl2axi4_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(tl2axi4_auto_out_ar_bits_user),
    .auto_out_r_ready(tl2axi4_auto_out_r_ready),
    .auto_out_r_valid(tl2axi4_auto_out_r_valid),
    .auto_out_r_bits_id(tl2axi4_auto_out_r_bits_id),
    .auto_out_r_bits_data(tl2axi4_auto_out_r_bits_data),
    .auto_out_r_bits_resp(tl2axi4_auto_out_r_bits_resp),
    .auto_out_r_bits_user(tl2axi4_auto_out_r_bits_user),
    .auto_out_r_bits_last(tl2axi4_auto_out_r_bits_last)
  );
  TLBuffer_16 buffer ( // @[Buffer.scala 69:28:boom.system.TestHarness.MegaBoomConfig.fir@31761.4]
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
  );
  assign auto_buffer_in_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_buffer_in_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_buffer_in_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_buffer_in_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_buffer_in_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_buffer_in_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_buffer_in_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_buffer_in_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_buffer_in_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign auto_axi4yank_out_aw_valid = axi4yank_auto_out_aw_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_id = axi4yank_auto_out_aw_bits_id; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_addr = axi4yank_auto_out_aw_bits_addr; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_len = axi4yank_auto_out_aw_bits_len; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_size = axi4yank_auto_out_aw_bits_size; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_burst = axi4yank_auto_out_aw_bits_burst; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_lock = axi4yank_auto_out_aw_bits_lock; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_cache = axi4yank_auto_out_aw_bits_cache; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_prot = axi4yank_auto_out_aw_bits_prot; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_aw_bits_qos = axi4yank_auto_out_aw_bits_qos; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_w_valid = axi4yank_auto_out_w_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_w_bits_data = axi4yank_auto_out_w_bits_data; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_w_bits_strb = axi4yank_auto_out_w_bits_strb; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_w_bits_last = axi4yank_auto_out_w_bits_last; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_b_ready = axi4yank_auto_out_b_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_valid = axi4yank_auto_out_ar_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_id = axi4yank_auto_out_ar_bits_id; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_addr = axi4yank_auto_out_ar_bits_addr; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_len = axi4yank_auto_out_ar_bits_len; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_size = axi4yank_auto_out_ar_bits_size; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_burst = axi4yank_auto_out_ar_bits_burst; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_lock = axi4yank_auto_out_ar_bits_lock; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_cache = axi4yank_auto_out_ar_bits_cache; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_prot = axi4yank_auto_out_ar_bits_prot; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_ar_bits_qos = axi4yank_auto_out_ar_bits_qos; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign auto_axi4yank_out_r_ready = axi4yank_auto_out_r_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@31747.4]
  assign axi4yank_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@31748.4]
  assign axi4yank_auto_in_aw_valid = axi4index_auto_out_aw_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_id = axi4index_auto_out_aw_bits_id; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_addr = axi4index_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_len = axi4index_auto_out_aw_bits_len; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_size = axi4index_auto_out_aw_bits_size; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_burst = axi4index_auto_out_aw_bits_burst; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_lock = axi4index_auto_out_aw_bits_lock; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_cache = axi4index_auto_out_aw_bits_cache; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_prot = axi4index_auto_out_aw_bits_prot; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_qos = axi4index_auto_out_aw_bits_qos; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_aw_bits_user = axi4index_auto_out_aw_bits_user; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_w_valid = axi4index_auto_out_w_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_w_bits_data = axi4index_auto_out_w_bits_data; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_w_bits_strb = axi4index_auto_out_w_bits_strb; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_w_bits_last = axi4index_auto_out_w_bits_last; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_b_ready = axi4index_auto_out_b_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_valid = axi4index_auto_out_ar_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_id = axi4index_auto_out_ar_bits_id; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_addr = axi4index_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_len = axi4index_auto_out_ar_bits_len; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_size = axi4index_auto_out_ar_bits_size; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_burst = axi4index_auto_out_ar_bits_burst; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_lock = axi4index_auto_out_ar_bits_lock; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_cache = axi4index_auto_out_ar_bits_cache; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_prot = axi4index_auto_out_ar_bits_prot; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_qos = axi4index_auto_out_ar_bits_qos; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_ar_bits_user = axi4index_auto_out_ar_bits_user; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_in_r_ready = axi4index_auto_out_r_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4yank_auto_out_aw_ready = auto_axi4yank_out_aw_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_w_ready = auto_axi4yank_out_w_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_b_valid = auto_axi4yank_out_b_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_b_bits_id = auto_axi4yank_out_b_bits_id; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_b_bits_resp = auto_axi4yank_out_b_bits_resp; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_ar_ready = auto_axi4yank_out_ar_ready; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_r_valid = auto_axi4yank_out_r_valid; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_r_bits_id = auto_axi4yank_out_r_bits_id; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_r_bits_data = auto_axi4yank_out_r_bits_data; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_r_bits_resp = auto_axi4yank_out_r_bits_resp; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4yank_auto_out_r_bits_last = auto_axi4yank_out_r_bits_last; // @[LazyModule.scala 173:49:boom.system.TestHarness.MegaBoomConfig.fir@31770.4]
  assign axi4index_auto_in_aw_valid = tl2axi4_auto_out_aw_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_id = tl2axi4_auto_out_aw_bits_id; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_addr = tl2axi4_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_len = tl2axi4_auto_out_aw_bits_len; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_size = tl2axi4_auto_out_aw_bits_size; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_burst = tl2axi4_auto_out_aw_bits_burst; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_lock = tl2axi4_auto_out_aw_bits_lock; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_cache = tl2axi4_auto_out_aw_bits_cache; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_prot = tl2axi4_auto_out_aw_bits_prot; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_qos = tl2axi4_auto_out_aw_bits_qos; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_aw_bits_user = tl2axi4_auto_out_aw_bits_user; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_w_valid = tl2axi4_auto_out_w_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_w_bits_data = tl2axi4_auto_out_w_bits_data; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_w_bits_strb = tl2axi4_auto_out_w_bits_strb; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_w_bits_last = tl2axi4_auto_out_w_bits_last; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_b_ready = tl2axi4_auto_out_b_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_valid = tl2axi4_auto_out_ar_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_id = tl2axi4_auto_out_ar_bits_id; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_addr = tl2axi4_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_len = tl2axi4_auto_out_ar_bits_len; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_size = tl2axi4_auto_out_ar_bits_size; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_burst = tl2axi4_auto_out_ar_bits_burst; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_lock = tl2axi4_auto_out_ar_bits_lock; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_cache = tl2axi4_auto_out_ar_bits_cache; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_prot = tl2axi4_auto_out_ar_bits_prot; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_qos = tl2axi4_auto_out_ar_bits_qos; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_ar_bits_user = tl2axi4_auto_out_ar_bits_user; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_in_r_ready = tl2axi4_auto_out_r_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign axi4index_auto_out_aw_ready = axi4yank_auto_in_aw_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_w_ready = axi4yank_auto_in_w_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_b_valid = axi4yank_auto_in_b_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_b_bits_id = axi4yank_auto_in_b_bits_id; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_b_bits_resp = axi4yank_auto_in_b_bits_resp; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_b_bits_user = axi4yank_auto_in_b_bits_user; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_ar_ready = axi4yank_auto_in_ar_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_r_valid = axi4yank_auto_in_r_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_r_bits_id = axi4yank_auto_in_r_bits_id; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_r_bits_data = axi4yank_auto_in_r_bits_data; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_r_bits_resp = axi4yank_auto_in_r_bits_resp; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_r_bits_user = axi4yank_auto_in_r_bits_user; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign axi4index_auto_out_r_bits_last = axi4yank_auto_in_r_bits_last; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31767.4]
  assign tl2axi4_clock = clock; // @[:boom.system.TestHarness.MegaBoomConfig.fir@31759.4]
  assign tl2axi4_reset = reset; // @[:boom.system.TestHarness.MegaBoomConfig.fir@31760.4]
  assign tl2axi4_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign tl2axi4_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign tl2axi4_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign tl2axi4_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign tl2axi4_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign tl2axi4_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign tl2axi4_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign tl2axi4_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign tl2axi4_auto_out_aw_ready = axi4index_auto_in_aw_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_w_ready = axi4index_auto_in_w_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_b_valid = axi4index_auto_in_b_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_b_bits_id = axi4index_auto_in_b_bits_id; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_b_bits_resp = axi4index_auto_in_b_bits_resp; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_b_bits_user = axi4index_auto_in_b_bits_user; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_ar_ready = axi4index_auto_in_ar_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_r_valid = axi4index_auto_in_r_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_r_bits_id = axi4index_auto_in_r_bits_id; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_r_bits_data = axi4index_auto_in_r_bits_data; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_r_bits_resp = axi4index_auto_in_r_bits_resp; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_r_bits_user = axi4index_auto_in_r_bits_user; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign tl2axi4_auto_out_r_bits_last = axi4index_auto_in_r_bits_last; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31768.4]
  assign buffer_auto_in_a_valid = auto_buffer_in_a_valid; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign buffer_auto_in_a_bits_opcode = auto_buffer_in_a_bits_opcode; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign buffer_auto_in_a_bits_size = auto_buffer_in_a_bits_size; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign buffer_auto_in_a_bits_source = auto_buffer_in_a_bits_source; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign buffer_auto_in_a_bits_address = auto_buffer_in_a_bits_address; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign buffer_auto_in_a_bits_mask = auto_buffer_in_a_bits_mask; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign buffer_auto_in_a_bits_data = auto_buffer_in_a_bits_data; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign buffer_auto_in_d_ready = auto_buffer_in_d_ready; // @[LazyModule.scala 173:31:boom.system.TestHarness.MegaBoomConfig.fir@31771.4]
  assign buffer_auto_out_a_ready = tl2axi4_auto_in_a_ready; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign buffer_auto_out_d_valid = tl2axi4_auto_in_d_valid; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign buffer_auto_out_d_bits_opcode = tl2axi4_auto_in_d_bits_opcode; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign buffer_auto_out_d_bits_param = 2'h0; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign buffer_auto_out_d_bits_size = tl2axi4_auto_in_d_bits_size; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign buffer_auto_out_d_bits_source = tl2axi4_auto_in_d_bits_source; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign buffer_auto_out_d_bits_denied = tl2axi4_auto_in_d_bits_denied; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign buffer_auto_out_d_bits_data = tl2axi4_auto_in_d_bits_data; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
  assign buffer_auto_out_d_bits_corrupt = tl2axi4_auto_in_d_bits_corrupt; // @[LazyModule.scala 167:31:boom.system.TestHarness.MegaBoomConfig.fir@31769.4]
endmodule
