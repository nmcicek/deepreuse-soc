module TLBuffer_33( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291938.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291939.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291940.4]
  output        auto_in_a_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input         auto_in_a_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [2:0]  auto_in_a_bits_opcode, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [2:0]  auto_in_a_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [6:0]  auto_in_a_bits_source, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [31:0] auto_in_a_bits_address, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [7:0]  auto_in_a_bits_mask, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [63:0] auto_in_a_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input         auto_in_d_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output        auto_in_d_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [2:0]  auto_in_d_bits_opcode, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [1:0]  auto_in_d_bits_param, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [2:0]  auto_in_d_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [6:0]  auto_in_d_bits_source, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output        auto_in_d_bits_denied, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [63:0] auto_in_d_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output        auto_in_d_bits_corrupt, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input         auto_out_a_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output        auto_out_a_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [2:0]  auto_out_a_bits_opcode, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [2:0]  auto_out_a_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [6:0]  auto_out_a_bits_source, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [31:0] auto_out_a_bits_address, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [7:0]  auto_out_a_bits_mask, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output [63:0] auto_out_a_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  output        auto_out_d_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input         auto_out_d_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [2:0]  auto_out_d_bits_opcode, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [2:0]  auto_out_d_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [6:0]  auto_out_d_bits_source, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input         auto_out_d_bits_denied, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input  [63:0] auto_out_d_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
  input         auto_out_d_bits_corrupt // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291941.4]
);
  wire  Queue_clock; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire  Queue_reset; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [2:0] Queue_io_enq_bits_opcode; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [2:0] Queue_io_enq_bits_size; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [6:0] Queue_io_enq_bits_source; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [31:0] Queue_io_enq_bits_address; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [7:0] Queue_io_enq_bits_mask; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [63:0] Queue_io_enq_bits_data; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [2:0] Queue_io_deq_bits_opcode; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [2:0] Queue_io_deq_bits_size; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [6:0] Queue_io_deq_bits_source; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [31:0] Queue_io_deq_bits_address; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [7:0] Queue_io_deq_bits_mask; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire [63:0] Queue_io_deq_bits_data; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
  wire  Queue_1_clock; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_reset; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [2:0] Queue_1_io_enq_bits_opcode; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [2:0] Queue_1_io_enq_bits_size; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [6:0] Queue_1_io_enq_bits_source; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_io_enq_bits_denied; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [63:0] Queue_1_io_enq_bits_data; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_io_enq_bits_corrupt; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [2:0] Queue_1_io_deq_bits_opcode; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [1:0] Queue_1_io_deq_bits_param; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [2:0] Queue_1_io_deq_bits_size; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [6:0] Queue_1_io_deq_bits_source; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_io_deq_bits_denied; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire [63:0] Queue_1_io_deq_bits_data; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  wire  Queue_1_io_deq_bits_corrupt; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
  Queue_42 Queue ( // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291952.4]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data)
  );
  Queue_43 Queue_1 ( // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291966.4]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_denied(Queue_1_io_enq_bits_denied),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_corrupt(Queue_1_io_enq_bits_corrupt),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_1_io_deq_bits_param),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_denied(Queue_1_io_deq_bits_denied),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_corrupt(Queue_1_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_in_d_valid = Queue_1_io_deq_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_in_d_bits_opcode = Queue_1_io_deq_bits_opcode; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_in_d_bits_param = Queue_1_io_deq_bits_param; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_in_d_bits_size = Queue_1_io_deq_bits_size; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_in_d_bits_source = Queue_1_io_deq_bits_source; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_in_d_bits_denied = Queue_1_io_deq_bits_denied; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_in_d_bits_data = Queue_1_io_deq_bits_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_in_d_bits_corrupt = Queue_1_io_deq_bits_corrupt; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291951.4]
  assign auto_out_a_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291950.4]
  assign auto_out_a_bits_opcode = Queue_io_deq_bits_opcode; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291950.4]
  assign auto_out_a_bits_size = Queue_io_deq_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291950.4]
  assign auto_out_a_bits_source = Queue_io_deq_bits_source; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291950.4]
  assign auto_out_a_bits_address = Queue_io_deq_bits_address; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291950.4]
  assign auto_out_a_bits_mask = Queue_io_deq_bits_mask; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291950.4]
  assign auto_out_a_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291950.4]
  assign auto_out_d_ready = Queue_1_io_enq_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291950.4]
  assign Queue_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291953.4]
  assign Queue_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291954.4]
  assign Queue_io_enq_valid = auto_in_a_valid; // @[Decoupled.scala 294:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291955.4]
  assign Queue_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291963.4]
  assign Queue_io_enq_bits_size = auto_in_a_bits_size; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291961.4]
  assign Queue_io_enq_bits_source = auto_in_a_bits_source; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291960.4]
  assign Queue_io_enq_bits_address = auto_in_a_bits_address; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291959.4]
  assign Queue_io_enq_bits_mask = auto_in_a_bits_mask; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291958.4]
  assign Queue_io_enq_bits_data = auto_in_a_bits_data; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291957.4]
  assign Queue_io_deq_ready = auto_out_a_ready; // @[Buffer.scala 38:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291965.4]
  assign Queue_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291967.4]
  assign Queue_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291968.4]
  assign Queue_1_io_enq_valid = auto_out_d_valid; // @[Decoupled.scala 294:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291969.4]
  assign Queue_1_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291977.4]
  assign Queue_1_io_enq_bits_size = auto_out_d_bits_size; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291975.4]
  assign Queue_1_io_enq_bits_source = auto_out_d_bits_source; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291974.4]
  assign Queue_1_io_enq_bits_denied = auto_out_d_bits_denied; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291972.4]
  assign Queue_1_io_enq_bits_data = auto_out_d_bits_data; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291971.4]
  assign Queue_1_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291970.4]
  assign Queue_1_io_deq_ready = auto_in_d_ready; // @[Buffer.scala 39:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291979.4]
endmodule
module Queue_44( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291987.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291988.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291989.4]
  output        io_enq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  input         io_enq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  input  [63:0] io_enq_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  input  [7:0]  io_enq_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  input         io_enq_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  input         io_deq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  output        io_deq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  output [63:0] io_deq_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  output [7:0]  io_deq_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
  output        io_deq_bits_last // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291990.4]
);
  reg [63:0] _T_35_data [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  reg [63:0] _RAND_0;
  wire [63:0] _T_35_data__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_data__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire [63:0] _T_35_data__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_data__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_data__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_data__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  reg [7:0] _T_35_strb [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  reg [31:0] _RAND_1;
  wire [7:0] _T_35_strb__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_strb__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire [7:0] _T_35_strb__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_strb__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_strb__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_strb__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  reg  _T_35_last [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  reg [31:0] _RAND_2;
  wire  _T_35_last__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_last__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_last__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_last__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_last__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  wire  _T_35_last__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  reg  _T_37; // @[Decoupled.scala 217:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291993.4]
  reg [31:0] _RAND_3;
  wire  _T_39; // @[Decoupled.scala 220:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291995.4]
  wire  _T_42; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291998.4]
  wire  _T_45; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292001.4]
  wire  _GEN_9; // @[Decoupled.scala 245:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292032.6]
  wire  _GEN_14; // @[Decoupled.scala 242:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292027.4]
  wire  _GEN_13; // @[Decoupled.scala 242:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292027.4]
  wire  _T_49; // @[Decoupled.scala 232:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292012.4]
  wire  _T_50; // @[Decoupled.scala 236:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292016.4]
  assign _T_35_data__T_52_addr = 1'h0;
  assign _T_35_data__T_52_data = _T_35_data[_T_35_data__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  assign _T_35_data__T_48_data = io_enq_bits_data;
  assign _T_35_data__T_48_addr = 1'h0;
  assign _T_35_data__T_48_mask = 1'h1;
  assign _T_35_data__T_48_en = _T_39 ? _GEN_9 : _T_42;
  assign _T_35_strb__T_52_addr = 1'h0;
  assign _T_35_strb__T_52_data = _T_35_strb[_T_35_strb__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  assign _T_35_strb__T_48_data = io_enq_bits_strb;
  assign _T_35_strb__T_48_addr = 1'h0;
  assign _T_35_strb__T_48_mask = 1'h1;
  assign _T_35_strb__T_48_en = _T_39 ? _GEN_9 : _T_42;
  assign _T_35_last__T_52_addr = 1'h0;
  assign _T_35_last__T_52_data = _T_35_last[_T_35_last__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
  assign _T_35_last__T_48_data = io_enq_bits_last;
  assign _T_35_last__T_48_addr = 1'h0;
  assign _T_35_last__T_48_mask = 1'h1;
  assign _T_35_last__T_48_en = _T_39 ? _GEN_9 : _T_42;
  assign _T_39 = _T_37 == 1'h0; // @[Decoupled.scala 220:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291995.4]
  assign _T_42 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291998.4]
  assign _T_45 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292001.4]
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_42; // @[Decoupled.scala 245:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292032.6]
  assign _GEN_14 = _T_39 ? _GEN_9 : _T_42; // @[Decoupled.scala 242:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292027.4]
  assign _GEN_13 = _T_39 ? 1'h0 : _T_45; // @[Decoupled.scala 242:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292027.4]
  assign _T_49 = _GEN_14 != _GEN_13; // @[Decoupled.scala 232:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292012.4]
  assign _T_50 = _T_39 == 1'h0; // @[Decoupled.scala 236:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292016.4]
  assign io_enq_ready = _T_37 == 1'h0; // @[Decoupled.scala 237:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292019.4]
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_50; // @[Decoupled.scala 236:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292017.4 Decoupled.scala 241:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292025.6]
  assign io_deq_bits_data = _T_39 ? io_enq_bits_data : _T_35_data__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292023.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292030.6]
  assign io_deq_bits_strb = _T_39 ? io_enq_bits_strb : _T_35_strb__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292022.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292029.6]
  assign io_deq_bits_last = _T_39 ? io_enq_bits_last : _T_35_last__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292021.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292028.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_strb[initvar] = _RAND_1[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_37 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35_data__T_48_en & _T_35_data__T_48_mask) begin
      _T_35_data[_T_35_data__T_48_addr] <= _T_35_data__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
    end
    if(_T_35_strb__T_48_en & _T_35_strb__T_48_mask) begin
      _T_35_strb[_T_35_strb__T_48_addr] <= _T_35_strb__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
    end
    if(_T_35_last__T_48_en & _T_35_last__T_48_mask) begin
      _T_35_last[_T_35_last__T_48_addr] <= _T_35_last__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@291992.4]
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_49) begin
        if (_T_39) begin
          if (io_deq_ready) begin
            _T_37 <= 1'h0;
          end else begin
            _T_37 <= _T_42;
          end
        end else begin
          _T_37 <= _T_42;
        end
      end
    end
  end
endmodule
module Queue_45( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292043.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292044.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292045.4]
  output        io_enq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  input         io_enq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  input  [5:0]  io_enq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  input  [31:0] io_enq_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  input  [7:0]  io_enq_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  input  [2:0]  io_enq_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  input  [10:0] io_enq_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  input         io_enq_bits_wen, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  input         io_deq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output        io_deq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [5:0]  io_deq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [31:0] io_deq_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [7:0]  io_deq_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [2:0]  io_deq_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [1:0]  io_deq_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output        io_deq_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [3:0]  io_deq_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [2:0]  io_deq_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [3:0]  io_deq_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output [10:0] io_deq_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
  output        io_deq_bits_wen // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292046.4]
);
  reg [5:0] _T_35_id [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_0;
  wire [5:0] _T_35_id__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_id__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [5:0] _T_35_id__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_id__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_id__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_id__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _T_35_addr [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_1;
  wire [31:0] _T_35_addr__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_addr__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [31:0] _T_35_addr__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_addr__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_addr__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_addr__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [7:0] _T_35_len [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_2;
  wire [7:0] _T_35_len__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_len__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [7:0] _T_35_len__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_len__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_len__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_len__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [2:0] _T_35_size [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_3;
  wire [2:0] _T_35_size__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_size__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [2:0] _T_35_size__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_size__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_size__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_size__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [1:0] _T_35_burst [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_4;
  wire [1:0] _T_35_burst__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_burst__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [1:0] _T_35_burst__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_burst__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_burst__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_burst__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg  _T_35_lock [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_5;
  wire  _T_35_lock__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_lock__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_lock__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_lock__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_lock__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_lock__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [3:0] _T_35_cache [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_6;
  wire [3:0] _T_35_cache__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_cache__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [3:0] _T_35_cache__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_cache__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_cache__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_cache__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [2:0] _T_35_prot [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_7;
  wire [2:0] _T_35_prot__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_prot__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [2:0] _T_35_prot__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_prot__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_prot__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_prot__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [3:0] _T_35_qos [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_8;
  wire [3:0] _T_35_qos__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_qos__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [3:0] _T_35_qos__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_qos__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_qos__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_qos__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [10:0] _T_35_user [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_9;
  wire [10:0] _T_35_user__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_user__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire [10:0] _T_35_user__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_user__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_user__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_user__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg  _T_35_wen [0:0]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg [31:0] _RAND_10;
  wire  _T_35_wen__T_52_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_wen__T_52_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_wen__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_wen__T_48_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_wen__T_48_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  wire  _T_35_wen__T_48_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  reg  _T_37; // @[Decoupled.scala 217:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292049.4]
  reg [31:0] _RAND_11;
  wire  _T_39; // @[Decoupled.scala 220:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292051.4]
  wire  _T_42; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292054.4]
  wire  _T_45; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292057.4]
  wire  _GEN_17; // @[Decoupled.scala 245:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292112.6]
  wire  _GEN_30; // @[Decoupled.scala 242:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292099.4]
  wire  _GEN_29; // @[Decoupled.scala 242:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292099.4]
  wire  _T_49; // @[Decoupled.scala 232:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292076.4]
  wire  _T_50; // @[Decoupled.scala 236:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292080.4]
  assign _T_35_id__T_52_addr = 1'h0;
  assign _T_35_id__T_52_data = _T_35_id[_T_35_id__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_id__T_48_data = io_enq_bits_id;
  assign _T_35_id__T_48_addr = 1'h0;
  assign _T_35_id__T_48_mask = 1'h1;
  assign _T_35_id__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_addr__T_52_addr = 1'h0;
  assign _T_35_addr__T_52_data = _T_35_addr[_T_35_addr__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_addr__T_48_data = io_enq_bits_addr;
  assign _T_35_addr__T_48_addr = 1'h0;
  assign _T_35_addr__T_48_mask = 1'h1;
  assign _T_35_addr__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_len__T_52_addr = 1'h0;
  assign _T_35_len__T_52_data = _T_35_len[_T_35_len__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_len__T_48_data = io_enq_bits_len;
  assign _T_35_len__T_48_addr = 1'h0;
  assign _T_35_len__T_48_mask = 1'h1;
  assign _T_35_len__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_size__T_52_addr = 1'h0;
  assign _T_35_size__T_52_data = _T_35_size[_T_35_size__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_size__T_48_data = io_enq_bits_size;
  assign _T_35_size__T_48_addr = 1'h0;
  assign _T_35_size__T_48_mask = 1'h1;
  assign _T_35_size__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_burst__T_52_addr = 1'h0;
  assign _T_35_burst__T_52_data = _T_35_burst[_T_35_burst__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_burst__T_48_data = 2'h1;
  assign _T_35_burst__T_48_addr = 1'h0;
  assign _T_35_burst__T_48_mask = 1'h1;
  assign _T_35_burst__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_lock__T_52_addr = 1'h0;
  assign _T_35_lock__T_52_data = _T_35_lock[_T_35_lock__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_lock__T_48_data = 1'h0;
  assign _T_35_lock__T_48_addr = 1'h0;
  assign _T_35_lock__T_48_mask = 1'h1;
  assign _T_35_lock__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_cache__T_52_addr = 1'h0;
  assign _T_35_cache__T_52_data = _T_35_cache[_T_35_cache__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_cache__T_48_data = 4'h0;
  assign _T_35_cache__T_48_addr = 1'h0;
  assign _T_35_cache__T_48_mask = 1'h1;
  assign _T_35_cache__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_prot__T_52_addr = 1'h0;
  assign _T_35_prot__T_52_data = _T_35_prot[_T_35_prot__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_prot__T_48_data = 3'h1;
  assign _T_35_prot__T_48_addr = 1'h0;
  assign _T_35_prot__T_48_mask = 1'h1;
  assign _T_35_prot__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_qos__T_52_addr = 1'h0;
  assign _T_35_qos__T_52_data = _T_35_qos[_T_35_qos__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_qos__T_48_data = 4'h0;
  assign _T_35_qos__T_48_addr = 1'h0;
  assign _T_35_qos__T_48_mask = 1'h1;
  assign _T_35_qos__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_user__T_52_addr = 1'h0;
  assign _T_35_user__T_52_data = _T_35_user[_T_35_user__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_user__T_48_data = io_enq_bits_user;
  assign _T_35_user__T_48_addr = 1'h0;
  assign _T_35_user__T_48_mask = 1'h1;
  assign _T_35_user__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_35_wen__T_52_addr = 1'h0;
  assign _T_35_wen__T_52_data = _T_35_wen[_T_35_wen__T_52_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
  assign _T_35_wen__T_48_data = io_enq_bits_wen;
  assign _T_35_wen__T_48_addr = 1'h0;
  assign _T_35_wen__T_48_mask = 1'h1;
  assign _T_35_wen__T_48_en = _T_39 ? _GEN_17 : _T_42;
  assign _T_39 = _T_37 == 1'h0; // @[Decoupled.scala 220:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292051.4]
  assign _T_42 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292054.4]
  assign _T_45 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292057.4]
  assign _GEN_17 = io_deq_ready ? 1'h0 : _T_42; // @[Decoupled.scala 245:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292112.6]
  assign _GEN_30 = _T_39 ? _GEN_17 : _T_42; // @[Decoupled.scala 242:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292099.4]
  assign _GEN_29 = _T_39 ? 1'h0 : _T_45; // @[Decoupled.scala 242:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292099.4]
  assign _T_49 = _GEN_30 != _GEN_29; // @[Decoupled.scala 232:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292076.4]
  assign _T_50 = _T_39 == 1'h0; // @[Decoupled.scala 236:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292080.4]
  assign io_enq_ready = _T_37 == 1'h0; // @[Decoupled.scala 237:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292083.4]
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_50; // @[Decoupled.scala 236:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292081.4 Decoupled.scala 241:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292097.6]
  assign io_deq_bits_id = _T_39 ? io_enq_bits_id : _T_35_id__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292095.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292110.6]
  assign io_deq_bits_addr = _T_39 ? io_enq_bits_addr : _T_35_addr__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292094.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292109.6]
  assign io_deq_bits_len = _T_39 ? io_enq_bits_len : _T_35_len__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292093.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292108.6]
  assign io_deq_bits_size = _T_39 ? io_enq_bits_size : _T_35_size__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292092.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292107.6]
  assign io_deq_bits_burst = _T_39 ? 2'h1 : _T_35_burst__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292091.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292106.6]
  assign io_deq_bits_lock = _T_39 ? 1'h0 : _T_35_lock__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292090.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292105.6]
  assign io_deq_bits_cache = _T_39 ? 4'h0 : _T_35_cache__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292089.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292104.6]
  assign io_deq_bits_prot = _T_39 ? 3'h1 : _T_35_prot__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292088.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292103.6]
  assign io_deq_bits_qos = _T_39 ? 4'h0 : _T_35_qos__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292087.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292102.6]
  assign io_deq_bits_user = _T_39 ? io_enq_bits_user : _T_35_user__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292086.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292101.6]
  assign io_deq_bits_wen = _T_39 ? io_enq_bits_wen : _T_35_wen__T_52_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292085.4 Decoupled.scala 243:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292100.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_id[initvar] = _RAND_0[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_addr[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_user[initvar] = _RAND_9[10:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_35_wen[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_37 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35_id__T_48_en & _T_35_id__T_48_mask) begin
      _T_35_id[_T_35_id__T_48_addr] <= _T_35_id__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_addr__T_48_en & _T_35_addr__T_48_mask) begin
      _T_35_addr[_T_35_addr__T_48_addr] <= _T_35_addr__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_len__T_48_en & _T_35_len__T_48_mask) begin
      _T_35_len[_T_35_len__T_48_addr] <= _T_35_len__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_size__T_48_en & _T_35_size__T_48_mask) begin
      _T_35_size[_T_35_size__T_48_addr] <= _T_35_size__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_burst__T_48_en & _T_35_burst__T_48_mask) begin
      _T_35_burst[_T_35_burst__T_48_addr] <= _T_35_burst__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_lock__T_48_en & _T_35_lock__T_48_mask) begin
      _T_35_lock[_T_35_lock__T_48_addr] <= _T_35_lock__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_cache__T_48_en & _T_35_cache__T_48_mask) begin
      _T_35_cache[_T_35_cache__T_48_addr] <= _T_35_cache__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_prot__T_48_en & _T_35_prot__T_48_mask) begin
      _T_35_prot[_T_35_prot__T_48_addr] <= _T_35_prot__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_qos__T_48_en & _T_35_qos__T_48_mask) begin
      _T_35_qos[_T_35_qos__T_48_addr] <= _T_35_qos__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_user__T_48_en & _T_35_user__T_48_mask) begin
      _T_35_user[_T_35_user__T_48_addr] <= _T_35_user__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if(_T_35_wen__T_48_en & _T_35_wen__T_48_mask) begin
      _T_35_wen[_T_35_wen__T_48_addr] <= _T_35_wen__T_48_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292048.4]
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_49) begin
        if (_T_39) begin
          if (io_deq_ready) begin
            _T_37 <= 1'h0;
          end else begin
            _T_37 <= _T_42;
          end
        end else begin
          _T_37 <= _T_42;
        end
      end
    end
  end
endmodule
module TLToAXI4( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292123.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292124.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292125.4]
  output        auto_in_a_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input         auto_in_a_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [2:0]  auto_in_a_bits_opcode, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [2:0]  auto_in_a_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [6:0]  auto_in_a_bits_source, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [31:0] auto_in_a_bits_address, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [7:0]  auto_in_a_bits_mask, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [63:0] auto_in_a_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input         auto_in_d_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_in_d_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [2:0]  auto_in_d_bits_opcode, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [2:0]  auto_in_d_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [6:0]  auto_in_d_bits_source, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_in_d_bits_denied, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [63:0] auto_in_d_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_in_d_bits_corrupt, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input         auto_out_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_out_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [5:0]  auto_out_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [31:0] auto_out_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [7:0]  auto_out_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [2:0]  auto_out_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_out_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [10:0] auto_out_aw_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input         auto_out_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_out_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [63:0] auto_out_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [7:0]  auto_out_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_out_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_out_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input         auto_out_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [5:0]  auto_out_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [10:0] auto_out_b_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input         auto_out_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_out_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [5:0]  auto_out_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [31:0] auto_out_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [7:0]  auto_out_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [2:0]  auto_out_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_out_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output [10:0] auto_out_ar_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  output        auto_out_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input         auto_out_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [5:0]  auto_out_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [63:0] auto_out_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input  [10:0] auto_out_r_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
  input         auto_out_r_bits_last // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292126.4]
);
  wire  Queue_clock; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire  Queue_reset; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire [63:0] Queue_io_enq_bits_data; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire [7:0] Queue_io_enq_bits_strb; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire [63:0] Queue_io_deq_bits_data; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire [7:0] Queue_io_deq_bits_strb; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
  wire  Queue_1_clock; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  Queue_1_reset; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [5:0] Queue_1_io_enq_bits_id; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [31:0] Queue_1_io_enq_bits_addr; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [7:0] Queue_1_io_enq_bits_len; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [2:0] Queue_1_io_enq_bits_size; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [10:0] Queue_1_io_enq_bits_user; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  Queue_1_io_enq_bits_wen; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [5:0] Queue_1_io_deq_bits_id; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [31:0] Queue_1_io_deq_bits_addr; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [7:0] Queue_1_io_deq_bits_len; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [2:0] Queue_1_io_deq_bits_size; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [1:0] Queue_1_io_deq_bits_burst; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  Queue_1_io_deq_bits_lock; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [3:0] Queue_1_io_deq_bits_cache; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [2:0] Queue_1_io_deq_bits_prot; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [3:0] Queue_1_io_deq_bits_qos; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire [10:0] Queue_1_io_deq_bits_user; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  Queue_1_io_deq_bits_wen; // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
  wire  _T_887; // @[Edges.scala 92:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292466.4]
  wire  _T_888; // @[Edges.scala 92:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292467.4]
  reg  _T_3099; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295452.4]
  reg [31:0] _RAND_0;
  reg  _T_3068; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295410.4]
  reg [31:0] _RAND_1;
  reg  _T_3037; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295368.4]
  reg [31:0] _RAND_2;
  reg  _T_3006; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295326.4]
  reg [31:0] _RAND_3;
  reg  _T_2975; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295284.4]
  reg [31:0] _RAND_4;
  reg  _T_2944; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295242.4]
  reg [31:0] _RAND_5;
  reg  _T_2913; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295200.4]
  reg [31:0] _RAND_6;
  reg  _T_2882; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295158.4]
  reg [31:0] _RAND_7;
  reg  _T_2851; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295116.4]
  reg [31:0] _RAND_8;
  reg  _T_2820; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295074.4]
  reg [31:0] _RAND_9;
  reg  _T_2789; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295032.4]
  reg [31:0] _RAND_10;
  reg  _T_2758; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294990.4]
  reg [31:0] _RAND_11;
  reg  _T_2727; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294948.4]
  reg [31:0] _RAND_12;
  reg  _T_2696; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294906.4]
  reg [31:0] _RAND_13;
  reg  _T_2665; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294864.4]
  reg [31:0] _RAND_14;
  reg  _T_2634; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294822.4]
  reg [31:0] _RAND_15;
  reg  _T_2603; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294780.4]
  reg [31:0] _RAND_16;
  reg  _T_2572; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294738.4]
  reg [31:0] _RAND_17;
  reg  _T_2541; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294696.4]
  reg [31:0] _RAND_18;
  reg  _T_2510; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294654.4]
  reg [31:0] _RAND_19;
  reg  _T_2479; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294612.4]
  reg [31:0] _RAND_20;
  reg  _T_2448; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294570.4]
  reg [31:0] _RAND_21;
  reg  _T_2417; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294528.4]
  reg [31:0] _RAND_22;
  reg  _T_2386; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294486.4]
  reg [31:0] _RAND_23;
  reg  _T_2355; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294444.4]
  reg [31:0] _RAND_24;
  reg  _T_2324; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294402.4]
  reg [31:0] _RAND_25;
  reg  _T_2293; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294360.4]
  reg [31:0] _RAND_26;
  reg  _T_2262; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294318.4]
  reg [31:0] _RAND_27;
  reg  _T_2231; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294276.4]
  reg [31:0] _RAND_28;
  reg  _T_2200; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294234.4]
  reg [31:0] _RAND_29;
  reg  _T_2169; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294192.4]
  reg [31:0] _RAND_30;
  reg  _T_2138; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294150.4]
  reg [31:0] _RAND_31;
  reg  _T_2107; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294108.4]
  reg [31:0] _RAND_32;
  reg  _T_2076; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294066.4]
  reg [31:0] _RAND_33;
  reg  _T_2045; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294024.4]
  reg [31:0] _RAND_34;
  reg  _T_2014; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293982.4]
  reg [31:0] _RAND_35;
  reg  _T_1983; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293940.4]
  reg [31:0] _RAND_36;
  reg  _T_1952; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293898.4]
  reg [31:0] _RAND_37;
  reg  _T_1921; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293856.4]
  reg [31:0] _RAND_38;
  reg  _T_1890; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293814.4]
  reg [31:0] _RAND_39;
  reg  _T_1859; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293772.4]
  reg [31:0] _RAND_40;
  reg  _T_1828; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293730.4]
  reg [31:0] _RAND_41;
  reg  _T_1797; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293688.4]
  reg [31:0] _RAND_42;
  reg  _T_1766; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293646.4]
  reg [31:0] _RAND_43;
  reg  _T_1735; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293604.4]
  reg [31:0] _RAND_44;
  reg  _T_1704; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293562.4]
  reg [31:0] _RAND_45;
  reg  _T_1673; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293520.4]
  reg [31:0] _RAND_46;
  reg  _T_1642; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293478.4]
  reg [31:0] _RAND_47;
  reg  _T_1611; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293436.4]
  reg [31:0] _RAND_48;
  reg  _T_1580; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293394.4]
  reg [31:0] _RAND_49;
  reg  _T_1549; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293352.4]
  reg [31:0] _RAND_50;
  reg  _T_1518; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293310.4]
  reg [31:0] _RAND_51;
  reg  _T_1487; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293268.4]
  reg [31:0] _RAND_52;
  reg  _T_1456; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293226.4]
  reg [31:0] _RAND_53;
  reg  _T_1425; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293184.4]
  reg [31:0] _RAND_54;
  reg  _T_1394; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293142.4]
  reg [31:0] _RAND_55;
  reg  _T_1363; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293100.4]
  reg [31:0] _RAND_56;
  reg  _T_1332; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293058.4]
  reg [31:0] _RAND_57;
  reg  _T_1301; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293016.4]
  reg [31:0] _RAND_58;
  reg  _T_1270; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292974.4]
  reg [31:0] _RAND_59;
  reg  _T_1239; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292932.4]
  reg [31:0] _RAND_60;
  reg  _T_1208; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292890.4]
  reg [31:0] _RAND_61;
  reg  _T_1177; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292848.4]
  reg [31:0] _RAND_62;
  reg  _T_1146; // @[ToAXI4.scala 225:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292806.4]
  reg [31:0] _RAND_63;
  wire  _GEN_132; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_133; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_134; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_135; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_136; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_137; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_138; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_139; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_140; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_141; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_142; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_143; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_144; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_145; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_146; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_147; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_148; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_149; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_150; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_151; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_152; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_153; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_154; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_155; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_156; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_157; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_158; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_159; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_160; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_161; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_162; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_163; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_164; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_165; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_166; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_167; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_168; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_169; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_170; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_171; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_172; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_173; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_174; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_175; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_176; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_177; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_178; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_179; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_180; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_181; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_182; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_183; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_184; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_185; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_186; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_187; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_188; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_189; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_190; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_191; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_192; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_193; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_194; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_195; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_196; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_197; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_198; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_199; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_200; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_201; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_202; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_203; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_204; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_205; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_206; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_207; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_208; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_209; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_210; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_211; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_212; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_213; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_214; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_215; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_216; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_217; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_218; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_219; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_220; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_221; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_222; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_223; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_224; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_225; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_226; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_227; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_228; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_229; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_230; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_231; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_232; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_233; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_234; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_235; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_236; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_237; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_238; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_239; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_240; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_241; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_242; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_243; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_244; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_245; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_246; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_247; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_248; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_249; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_250; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_251; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_252; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_253; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_254; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_255; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_256; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _GEN_257; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  reg [3:0] _T_899; // @[Edges.scala 229:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292477.4]
  reg [31:0] _RAND_64;
  wire  _T_903; // @[Edges.scala 231:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292481.4]
  wire  _T_969; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  wire  _T_970; // @[ToAXI4.scala 177:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292598.4]
  reg  _T_957; // @[ToAXI4.scala 160:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292573.4]
  reg [31:0] _RAND_65;
  wire  _T_930_ready; // @[ToAXI4.scala 146:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292515.4 Decoupled.scala 296:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292549.4]
  wire  _T_971; // @[ToAXI4.scala 177:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292599.4]
  wire  _T_933_ready; // @[ToAXI4.scala 147:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292517.4 Decoupled.scala 296:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292526.4]
  wire  _T_972; // @[ToAXI4.scala 177:70:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292600.4]
  wire  _T_973; // @[ToAXI4.scala 177:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292601.4]
  wire  _T_974; // @[ToAXI4.scala 177:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292602.4]
  wire  _T_889; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292468.4]
  wire [13:0] _T_891; // @[package.scala 185:77:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292470.4]
  wire [6:0] _T_892; // @[package.scala 185:82:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292471.4]
  wire [6:0] _T_893; // @[package.scala 185:46:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292472.4]
  wire [3:0] _T_894; // @[Edges.scala 220:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292473.4]
  wire [3:0] _T_897; // @[Edges.scala 221:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292476.4]
  wire [4:0] _T_900; // @[Edges.scala 230:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292478.4]
  wire [4:0] _T_901; // @[Edges.scala 230:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292479.4]
  wire [3:0] _T_902; // @[Edges.scala 230:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292480.4]
  wire  _T_904; // @[Edges.scala 232:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292482.4]
  wire  _T_905; // @[Edges.scala 232:47:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292483.4]
  wire  _T_906; // @[Edges.scala 232:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292484.4]
  wire [9:0] _GEN_325; // @[ToAXI4.scala 134:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292509.4]
  wire [9:0] _T_920; // @[ToAXI4.scala 134:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292509.4]
  wire [9:0] _GEN_326; // @[ToAXI4.scala 134:45:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292510.4]
  wire [9:0] _T_921; // @[ToAXI4.scala 134:45:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292510.4]
  wire [6:0] _T_922; // @[ToAXI4.scala 137:50:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292511.4]
  wire [2:0] _T_923; // @[ToAXI4.scala 138:50:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292512.4]
  wire [6:0] _T_924; // @[ToAXI4.scala 141:50:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292513.4]
  wire [2:0] _T_925; // @[ToAXI4.scala 142:50:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292514.4]
  wire  _T_948_bits_wen; // @[Decoupled.scala 314:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292550.4 Decoupled.scala 315:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292551.4]
  wire  _T_952; // @[ToAXI4.scala 154:42:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292566.4]
  wire  _T_948_valid; // @[Decoupled.scala 314:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292550.4 Decoupled.scala 316:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292562.4]
  wire  _T_959; // @[ToAXI4.scala 161:38:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292576.6]
  wire [5:0] _GEN_4; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_5; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_6; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_7; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_8; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_9; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_10; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_11; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_12; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_13; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_14; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_15; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_16; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_17; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_18; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_19; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_20; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_21; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_22; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_23; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_24; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_25; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_26; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_27; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_28; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_29; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_30; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_31; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_32; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_33; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_34; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_35; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_36; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_37; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_38; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_39; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_40; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_41; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_42; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_43; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_44; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_45; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_46; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_47; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_48; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_49; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_50; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_51; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_52; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_53; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_54; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_55; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_56; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_57; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_58; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_59; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_60; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_61; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_62; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_63; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_64; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_65; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_66; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_67; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_68; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_69; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_70; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_71; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_72; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_73; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_74; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_75; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_76; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_77; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_78; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_79; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_80; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_81; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_82; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_83; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_84; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_85; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_86; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_87; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_88; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_89; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_90; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_91; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_92; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_93; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_94; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_95; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_96; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_97; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_98; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_99; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_100; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_101; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_102; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_103; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_104; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_105; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_106; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_107; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_108; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_109; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_110; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_111; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_112; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_113; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_114; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_115; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_116; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_117; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_118; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_119; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_120; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_121; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_122; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_123; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_124; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_125; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_126; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_127; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_128; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [5:0] _GEN_129; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  wire [17:0] _T_962; // @[package.scala 185:77:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292583.4]
  wire [10:0] _T_963; // @[package.scala 185:82:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292584.4]
  wire [10:0] _T_964; // @[package.scala 185:46:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292585.4]
  wire  _T_966; // @[ToAXI4.scala 168:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292588.4]
  wire  _T_976; // @[ToAXI4.scala 178:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292605.4]
  wire  _T_977; // @[ToAXI4.scala 178:61:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292606.4]
  wire  _T_978; // @[ToAXI4.scala 178:69:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292607.4]
  wire  _T_979; // @[ToAXI4.scala 178:51:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292608.4]
  wire  _T_980; // @[ToAXI4.scala 178:45:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292609.4]
  wire  _T_983; // @[ToAXI4.scala 180:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292613.4]
  reg  _T_987; // @[ToAXI4.scala 187:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292620.4]
  reg [31:0] _RAND_66;
  wire  _T_988; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292621.4]
  wire  _T_989; // @[ToAXI4.scala 188:42:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292623.6]
  wire  _T_990; // @[ToAXI4.scala 190:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292626.4]
  wire  _T_991; // @[ToAXI4.scala 193:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292628.4]
  wire  _T_993; // @[ToAXI4.scala 194:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292631.4]
  reg  _T_995; // @[ToAXI4.scala 199:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292633.4]
  reg [31:0] _RAND_67;
  wire  _T_997; // @[ToAXI4.scala 201:39:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292638.4]
  reg  _T_999; // @[Reg.scala 11:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292639.4]
  reg [31:0] _RAND_68;
  wire  _GEN_260; // @[Reg.scala 12:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292640.4]
  wire  _T_1001; // @[ToAXI4.scala 202:39:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292644.4]
  wire  _T_1002; // @[ToAXI4.scala 203:39:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292645.4]
  wire  _T_1003; // @[ToAXI4.scala 205:100:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292646.4]
  wire [63:0] _T_1010; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292671.4]
  wire  _T_1012; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292673.4]
  wire  _T_1013; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292674.4]
  wire  _T_1014; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292675.4]
  wire  _T_1015; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292676.4]
  wire  _T_1016; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292677.4]
  wire  _T_1017; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292678.4]
  wire  _T_1018; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292679.4]
  wire  _T_1019; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292680.4]
  wire  _T_1020; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292681.4]
  wire  _T_1021; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292682.4]
  wire  _T_1022; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292683.4]
  wire  _T_1023; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292684.4]
  wire  _T_1024; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292685.4]
  wire  _T_1025; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292686.4]
  wire  _T_1026; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292687.4]
  wire  _T_1027; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292688.4]
  wire  _T_1028; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292689.4]
  wire  _T_1029; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292690.4]
  wire  _T_1030; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292691.4]
  wire  _T_1031; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292692.4]
  wire  _T_1032; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292693.4]
  wire  _T_1033; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292694.4]
  wire  _T_1034; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292695.4]
  wire  _T_1035; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292696.4]
  wire  _T_1036; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292697.4]
  wire  _T_1037; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292698.4]
  wire  _T_1038; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292699.4]
  wire  _T_1039; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292700.4]
  wire  _T_1040; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292701.4]
  wire  _T_1041; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292702.4]
  wire  _T_1042; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292703.4]
  wire  _T_1043; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292704.4]
  wire  _T_1044; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292705.4]
  wire  _T_1045; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292706.4]
  wire  _T_1046; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292707.4]
  wire  _T_1047; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292708.4]
  wire  _T_1048; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292709.4]
  wire  _T_1049; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292710.4]
  wire  _T_1050; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292711.4]
  wire  _T_1051; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292712.4]
  wire  _T_1052; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292713.4]
  wire  _T_1053; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292714.4]
  wire  _T_1054; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292715.4]
  wire  _T_1055; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292716.4]
  wire  _T_1056; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292717.4]
  wire  _T_1057; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292718.4]
  wire  _T_1058; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292719.4]
  wire  _T_1059; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292720.4]
  wire  _T_1060; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292721.4]
  wire  _T_1061; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292722.4]
  wire  _T_1062; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292723.4]
  wire  _T_1063; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292724.4]
  wire  _T_1064; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292725.4]
  wire  _T_1065; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292726.4]
  wire  _T_1066; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292727.4]
  wire  _T_1067; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292728.4]
  wire  _T_1068; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292729.4]
  wire  _T_1069; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292730.4]
  wire  _T_1070; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292731.4]
  wire  _T_1071; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292732.4]
  wire  _T_1072; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292733.4]
  wire  _T_1073; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292734.4]
  wire  _T_1074; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292735.4]
  wire  _T_1075; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292736.4]
  wire [5:0] _T_1076; // @[ToAXI4.scala 214:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292737.4]
  wire [63:0] _T_1078; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292739.4]
  wire  _T_1080; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292741.4]
  wire  _T_1081; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292742.4]
  wire  _T_1082; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292743.4]
  wire  _T_1083; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292744.4]
  wire  _T_1084; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292745.4]
  wire  _T_1085; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292746.4]
  wire  _T_1086; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292747.4]
  wire  _T_1087; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292748.4]
  wire  _T_1088; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292749.4]
  wire  _T_1089; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292750.4]
  wire  _T_1090; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292751.4]
  wire  _T_1091; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292752.4]
  wire  _T_1092; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292753.4]
  wire  _T_1093; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292754.4]
  wire  _T_1094; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292755.4]
  wire  _T_1095; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292756.4]
  wire  _T_1096; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292757.4]
  wire  _T_1097; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292758.4]
  wire  _T_1098; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292759.4]
  wire  _T_1099; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292760.4]
  wire  _T_1100; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292761.4]
  wire  _T_1101; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292762.4]
  wire  _T_1102; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292763.4]
  wire  _T_1103; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292764.4]
  wire  _T_1104; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292765.4]
  wire  _T_1105; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292766.4]
  wire  _T_1106; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292767.4]
  wire  _T_1107; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292768.4]
  wire  _T_1108; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292769.4]
  wire  _T_1109; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292770.4]
  wire  _T_1110; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292771.4]
  wire  _T_1111; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292772.4]
  wire  _T_1112; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292773.4]
  wire  _T_1113; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292774.4]
  wire  _T_1114; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292775.4]
  wire  _T_1115; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292776.4]
  wire  _T_1116; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292777.4]
  wire  _T_1117; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292778.4]
  wire  _T_1118; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292779.4]
  wire  _T_1119; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292780.4]
  wire  _T_1120; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292781.4]
  wire  _T_1121; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292782.4]
  wire  _T_1122; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292783.4]
  wire  _T_1123; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292784.4]
  wire  _T_1124; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292785.4]
  wire  _T_1125; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292786.4]
  wire  _T_1126; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292787.4]
  wire  _T_1127; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292788.4]
  wire  _T_1128; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292789.4]
  wire  _T_1129; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292790.4]
  wire  _T_1130; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292791.4]
  wire  _T_1131; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292792.4]
  wire  _T_1132; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292793.4]
  wire  _T_1133; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292794.4]
  wire  _T_1134; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292795.4]
  wire  _T_1135; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292796.4]
  wire  _T_1136; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292797.4]
  wire  _T_1137; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292798.4]
  wire  _T_1138; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292799.4]
  wire  _T_1139; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292800.4]
  wire  _T_1140; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292801.4]
  wire  _T_1141; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292802.4]
  wire  _T_1142; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292803.4]
  wire  _T_1143; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292804.4]
  wire  _T_1144; // @[ToAXI4.scala 215:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292805.4]
  wire  _T_1150; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292809.4]
  wire  _T_1151; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292810.4]
  wire  _T_1152; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292811.4]
  wire  _T_1153; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292812.4]
  wire  _T_1154; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292813.4]
  wire  _T_1156; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292815.4]
  wire [1:0] _T_1157; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292816.4]
  wire [1:0] _T_1158; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292817.4]
  wire  _T_1159; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292818.4]
  wire  _T_1160; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292820.4]
  wire  _T_1162; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292822.4]
  wire  _T_1164; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292824.4]
  wire  _T_1165; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292825.4]
  wire  _T_1166; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292830.4]
  wire  _T_1167; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292831.4]
  wire  _T_1168; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292832.4]
  wire  _T_1170; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292834.4]
  wire  _T_1171; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292835.4]
  wire  _T_1182; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292852.4]
  wire  _T_1183; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292853.4]
  wire  _T_1185; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292855.4]
  wire  _T_1187; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292857.4]
  wire [1:0] _T_1188; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292858.4]
  wire [1:0] _T_1189; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292859.4]
  wire  _T_1190; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292860.4]
  wire  _T_1191; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292862.4]
  wire  _T_1193; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292864.4]
  wire  _T_1195; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292866.4]
  wire  _T_1196; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292867.4]
  wire  _T_1197; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292872.4]
  wire  _T_1198; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292873.4]
  wire  _T_1199; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292874.4]
  wire  _T_1201; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292876.4]
  wire  _T_1202; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292877.4]
  wire  _T_1213; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292894.4]
  wire  _T_1214; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292895.4]
  wire  _T_1216; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292897.4]
  wire  _T_1218; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292899.4]
  wire [1:0] _T_1219; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292900.4]
  wire [1:0] _T_1220; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292901.4]
  wire  _T_1221; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292902.4]
  wire  _T_1222; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292904.4]
  wire  _T_1224; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292906.4]
  wire  _T_1226; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292908.4]
  wire  _T_1227; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292909.4]
  wire  _T_1228; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292914.4]
  wire  _T_1229; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292915.4]
  wire  _T_1230; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292916.4]
  wire  _T_1232; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292918.4]
  wire  _T_1233; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292919.4]
  wire  _T_1244; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292936.4]
  wire  _T_1245; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292937.4]
  wire  _T_1247; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292939.4]
  wire  _T_1249; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292941.4]
  wire [1:0] _T_1250; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292942.4]
  wire [1:0] _T_1251; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292943.4]
  wire  _T_1252; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292944.4]
  wire  _T_1253; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292946.4]
  wire  _T_1255; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292948.4]
  wire  _T_1257; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292950.4]
  wire  _T_1258; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292951.4]
  wire  _T_1259; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292956.4]
  wire  _T_1260; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292957.4]
  wire  _T_1261; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292958.4]
  wire  _T_1263; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292960.4]
  wire  _T_1264; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292961.4]
  wire  _T_1275; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292978.4]
  wire  _T_1276; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292979.4]
  wire  _T_1278; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292981.4]
  wire  _T_1280; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292983.4]
  wire [1:0] _T_1281; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292984.4]
  wire [1:0] _T_1282; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292985.4]
  wire  _T_1283; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292986.4]
  wire  _T_1284; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292988.4]
  wire  _T_1286; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292990.4]
  wire  _T_1288; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292992.4]
  wire  _T_1289; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292993.4]
  wire  _T_1290; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292998.4]
  wire  _T_1291; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292999.4]
  wire  _T_1292; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293000.4]
  wire  _T_1294; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293002.4]
  wire  _T_1295; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293003.4]
  wire  _T_1306; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293020.4]
  wire  _T_1307; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293021.4]
  wire  _T_1309; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293023.4]
  wire  _T_1311; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293025.4]
  wire [1:0] _T_1312; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293026.4]
  wire [1:0] _T_1313; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293027.4]
  wire  _T_1314; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293028.4]
  wire  _T_1315; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293030.4]
  wire  _T_1317; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293032.4]
  wire  _T_1319; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293034.4]
  wire  _T_1320; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293035.4]
  wire  _T_1321; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293040.4]
  wire  _T_1322; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293041.4]
  wire  _T_1323; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293042.4]
  wire  _T_1325; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293044.4]
  wire  _T_1326; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293045.4]
  wire  _T_1337; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293062.4]
  wire  _T_1338; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293063.4]
  wire  _T_1340; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293065.4]
  wire  _T_1342; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293067.4]
  wire [1:0] _T_1343; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293068.4]
  wire [1:0] _T_1344; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293069.4]
  wire  _T_1345; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293070.4]
  wire  _T_1346; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293072.4]
  wire  _T_1348; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293074.4]
  wire  _T_1350; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293076.4]
  wire  _T_1351; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293077.4]
  wire  _T_1352; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293082.4]
  wire  _T_1353; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293083.4]
  wire  _T_1354; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293084.4]
  wire  _T_1356; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293086.4]
  wire  _T_1357; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293087.4]
  wire  _T_1368; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293104.4]
  wire  _T_1369; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293105.4]
  wire  _T_1371; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293107.4]
  wire  _T_1373; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293109.4]
  wire [1:0] _T_1374; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293110.4]
  wire [1:0] _T_1375; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293111.4]
  wire  _T_1376; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293112.4]
  wire  _T_1377; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293114.4]
  wire  _T_1379; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293116.4]
  wire  _T_1381; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293118.4]
  wire  _T_1382; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293119.4]
  wire  _T_1383; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293124.4]
  wire  _T_1384; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293125.4]
  wire  _T_1385; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293126.4]
  wire  _T_1387; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293128.4]
  wire  _T_1388; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293129.4]
  wire  _T_1399; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293146.4]
  wire  _T_1400; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293147.4]
  wire  _T_1402; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293149.4]
  wire  _T_1404; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293151.4]
  wire [1:0] _T_1405; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293152.4]
  wire [1:0] _T_1406; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293153.4]
  wire  _T_1407; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293154.4]
  wire  _T_1408; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293156.4]
  wire  _T_1410; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293158.4]
  wire  _T_1412; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293160.4]
  wire  _T_1413; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293161.4]
  wire  _T_1414; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293166.4]
  wire  _T_1415; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293167.4]
  wire  _T_1416; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293168.4]
  wire  _T_1418; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293170.4]
  wire  _T_1419; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293171.4]
  wire  _T_1430; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293188.4]
  wire  _T_1431; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293189.4]
  wire  _T_1433; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293191.4]
  wire  _T_1435; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293193.4]
  wire [1:0] _T_1436; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293194.4]
  wire [1:0] _T_1437; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293195.4]
  wire  _T_1438; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293196.4]
  wire  _T_1439; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293198.4]
  wire  _T_1441; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293200.4]
  wire  _T_1443; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293202.4]
  wire  _T_1444; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293203.4]
  wire  _T_1445; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293208.4]
  wire  _T_1446; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293209.4]
  wire  _T_1447; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293210.4]
  wire  _T_1449; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293212.4]
  wire  _T_1450; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293213.4]
  wire  _T_1461; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293230.4]
  wire  _T_1462; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293231.4]
  wire  _T_1464; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293233.4]
  wire  _T_1466; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293235.4]
  wire [1:0] _T_1467; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293236.4]
  wire [1:0] _T_1468; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293237.4]
  wire  _T_1469; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293238.4]
  wire  _T_1470; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293240.4]
  wire  _T_1472; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293242.4]
  wire  _T_1474; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293244.4]
  wire  _T_1475; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293245.4]
  wire  _T_1476; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293250.4]
  wire  _T_1477; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293251.4]
  wire  _T_1478; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293252.4]
  wire  _T_1480; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293254.4]
  wire  _T_1481; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293255.4]
  wire  _T_1492; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293272.4]
  wire  _T_1493; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293273.4]
  wire  _T_1495; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293275.4]
  wire  _T_1497; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293277.4]
  wire [1:0] _T_1498; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293278.4]
  wire [1:0] _T_1499; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293279.4]
  wire  _T_1500; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293280.4]
  wire  _T_1501; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293282.4]
  wire  _T_1503; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293284.4]
  wire  _T_1505; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293286.4]
  wire  _T_1506; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293287.4]
  wire  _T_1507; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293292.4]
  wire  _T_1508; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293293.4]
  wire  _T_1509; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293294.4]
  wire  _T_1511; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293296.4]
  wire  _T_1512; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293297.4]
  wire  _T_1523; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293314.4]
  wire  _T_1524; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293315.4]
  wire  _T_1526; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293317.4]
  wire  _T_1528; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293319.4]
  wire [1:0] _T_1529; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293320.4]
  wire [1:0] _T_1530; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293321.4]
  wire  _T_1531; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293322.4]
  wire  _T_1532; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293324.4]
  wire  _T_1534; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293326.4]
  wire  _T_1536; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293328.4]
  wire  _T_1537; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293329.4]
  wire  _T_1538; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293334.4]
  wire  _T_1539; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293335.4]
  wire  _T_1540; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293336.4]
  wire  _T_1542; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293338.4]
  wire  _T_1543; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293339.4]
  wire  _T_1554; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293356.4]
  wire  _T_1555; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293357.4]
  wire  _T_1557; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293359.4]
  wire  _T_1559; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293361.4]
  wire [1:0] _T_1560; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293362.4]
  wire [1:0] _T_1561; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293363.4]
  wire  _T_1562; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293364.4]
  wire  _T_1563; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293366.4]
  wire  _T_1565; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293368.4]
  wire  _T_1567; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293370.4]
  wire  _T_1568; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293371.4]
  wire  _T_1569; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293376.4]
  wire  _T_1570; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293377.4]
  wire  _T_1571; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293378.4]
  wire  _T_1573; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293380.4]
  wire  _T_1574; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293381.4]
  wire  _T_1585; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293398.4]
  wire  _T_1586; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293399.4]
  wire  _T_1588; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293401.4]
  wire  _T_1590; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293403.4]
  wire [1:0] _T_1591; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293404.4]
  wire [1:0] _T_1592; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293405.4]
  wire  _T_1593; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293406.4]
  wire  _T_1594; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293408.4]
  wire  _T_1596; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293410.4]
  wire  _T_1598; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293412.4]
  wire  _T_1599; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293413.4]
  wire  _T_1600; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293418.4]
  wire  _T_1601; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293419.4]
  wire  _T_1602; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293420.4]
  wire  _T_1604; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293422.4]
  wire  _T_1605; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293423.4]
  wire  _T_1616; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293440.4]
  wire  _T_1617; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293441.4]
  wire  _T_1619; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293443.4]
  wire  _T_1621; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293445.4]
  wire [1:0] _T_1622; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293446.4]
  wire [1:0] _T_1623; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293447.4]
  wire  _T_1624; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293448.4]
  wire  _T_1625; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293450.4]
  wire  _T_1627; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293452.4]
  wire  _T_1629; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293454.4]
  wire  _T_1630; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293455.4]
  wire  _T_1631; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293460.4]
  wire  _T_1632; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293461.4]
  wire  _T_1633; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293462.4]
  wire  _T_1635; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293464.4]
  wire  _T_1636; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293465.4]
  wire  _T_1647; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293482.4]
  wire  _T_1648; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293483.4]
  wire  _T_1650; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293485.4]
  wire  _T_1652; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293487.4]
  wire [1:0] _T_1653; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293488.4]
  wire [1:0] _T_1654; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293489.4]
  wire  _T_1655; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293490.4]
  wire  _T_1656; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293492.4]
  wire  _T_1658; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293494.4]
  wire  _T_1660; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293496.4]
  wire  _T_1661; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293497.4]
  wire  _T_1662; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293502.4]
  wire  _T_1663; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293503.4]
  wire  _T_1664; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293504.4]
  wire  _T_1666; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293506.4]
  wire  _T_1667; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293507.4]
  wire  _T_1678; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293524.4]
  wire  _T_1679; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293525.4]
  wire  _T_1681; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293527.4]
  wire  _T_1683; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293529.4]
  wire [1:0] _T_1684; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293530.4]
  wire [1:0] _T_1685; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293531.4]
  wire  _T_1686; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293532.4]
  wire  _T_1687; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293534.4]
  wire  _T_1689; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293536.4]
  wire  _T_1691; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293538.4]
  wire  _T_1692; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293539.4]
  wire  _T_1693; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293544.4]
  wire  _T_1694; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293545.4]
  wire  _T_1695; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293546.4]
  wire  _T_1697; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293548.4]
  wire  _T_1698; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293549.4]
  wire  _T_1709; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293566.4]
  wire  _T_1710; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293567.4]
  wire  _T_1712; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293569.4]
  wire  _T_1714; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293571.4]
  wire [1:0] _T_1715; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293572.4]
  wire [1:0] _T_1716; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293573.4]
  wire  _T_1717; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293574.4]
  wire  _T_1718; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293576.4]
  wire  _T_1720; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293578.4]
  wire  _T_1722; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293580.4]
  wire  _T_1723; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293581.4]
  wire  _T_1724; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293586.4]
  wire  _T_1725; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293587.4]
  wire  _T_1726; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293588.4]
  wire  _T_1728; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293590.4]
  wire  _T_1729; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293591.4]
  wire  _T_1740; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293608.4]
  wire  _T_1741; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293609.4]
  wire  _T_1743; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293611.4]
  wire  _T_1745; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293613.4]
  wire [1:0] _T_1746; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293614.4]
  wire [1:0] _T_1747; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293615.4]
  wire  _T_1748; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293616.4]
  wire  _T_1749; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293618.4]
  wire  _T_1751; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293620.4]
  wire  _T_1753; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293622.4]
  wire  _T_1754; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293623.4]
  wire  _T_1755; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293628.4]
  wire  _T_1756; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293629.4]
  wire  _T_1757; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293630.4]
  wire  _T_1759; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293632.4]
  wire  _T_1760; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293633.4]
  wire  _T_1771; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293650.4]
  wire  _T_1772; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293651.4]
  wire  _T_1774; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293653.4]
  wire  _T_1776; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293655.4]
  wire [1:0] _T_1777; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293656.4]
  wire [1:0] _T_1778; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293657.4]
  wire  _T_1779; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293658.4]
  wire  _T_1780; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293660.4]
  wire  _T_1782; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293662.4]
  wire  _T_1784; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293664.4]
  wire  _T_1785; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293665.4]
  wire  _T_1786; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293670.4]
  wire  _T_1787; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293671.4]
  wire  _T_1788; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293672.4]
  wire  _T_1790; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293674.4]
  wire  _T_1791; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293675.4]
  wire  _T_1802; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293692.4]
  wire  _T_1803; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293693.4]
  wire  _T_1805; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293695.4]
  wire  _T_1807; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293697.4]
  wire [1:0] _T_1808; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293698.4]
  wire [1:0] _T_1809; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293699.4]
  wire  _T_1810; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293700.4]
  wire  _T_1811; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293702.4]
  wire  _T_1813; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293704.4]
  wire  _T_1815; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293706.4]
  wire  _T_1816; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293707.4]
  wire  _T_1817; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293712.4]
  wire  _T_1818; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293713.4]
  wire  _T_1819; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293714.4]
  wire  _T_1821; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293716.4]
  wire  _T_1822; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293717.4]
  wire  _T_1833; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293734.4]
  wire  _T_1834; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293735.4]
  wire  _T_1836; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293737.4]
  wire  _T_1838; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293739.4]
  wire [1:0] _T_1839; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293740.4]
  wire [1:0] _T_1840; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293741.4]
  wire  _T_1841; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293742.4]
  wire  _T_1842; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293744.4]
  wire  _T_1844; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293746.4]
  wire  _T_1846; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293748.4]
  wire  _T_1847; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293749.4]
  wire  _T_1848; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293754.4]
  wire  _T_1849; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293755.4]
  wire  _T_1850; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293756.4]
  wire  _T_1852; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293758.4]
  wire  _T_1853; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293759.4]
  wire  _T_1864; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293776.4]
  wire  _T_1865; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293777.4]
  wire  _T_1867; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293779.4]
  wire  _T_1869; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293781.4]
  wire [1:0] _T_1870; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293782.4]
  wire [1:0] _T_1871; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293783.4]
  wire  _T_1872; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293784.4]
  wire  _T_1873; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293786.4]
  wire  _T_1875; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293788.4]
  wire  _T_1877; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293790.4]
  wire  _T_1878; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293791.4]
  wire  _T_1879; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293796.4]
  wire  _T_1880; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293797.4]
  wire  _T_1881; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293798.4]
  wire  _T_1883; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293800.4]
  wire  _T_1884; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293801.4]
  wire  _T_1895; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293818.4]
  wire  _T_1896; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293819.4]
  wire  _T_1898; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293821.4]
  wire  _T_1900; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293823.4]
  wire [1:0] _T_1901; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293824.4]
  wire [1:0] _T_1902; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293825.4]
  wire  _T_1903; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293826.4]
  wire  _T_1904; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293828.4]
  wire  _T_1906; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293830.4]
  wire  _T_1908; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293832.4]
  wire  _T_1909; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293833.4]
  wire  _T_1910; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293838.4]
  wire  _T_1911; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293839.4]
  wire  _T_1912; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293840.4]
  wire  _T_1914; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293842.4]
  wire  _T_1915; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293843.4]
  wire  _T_1926; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293860.4]
  wire  _T_1927; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293861.4]
  wire  _T_1929; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293863.4]
  wire  _T_1931; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293865.4]
  wire [1:0] _T_1932; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293866.4]
  wire [1:0] _T_1933; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293867.4]
  wire  _T_1934; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293868.4]
  wire  _T_1935; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293870.4]
  wire  _T_1937; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293872.4]
  wire  _T_1939; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293874.4]
  wire  _T_1940; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293875.4]
  wire  _T_1941; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293880.4]
  wire  _T_1942; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293881.4]
  wire  _T_1943; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293882.4]
  wire  _T_1945; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293884.4]
  wire  _T_1946; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293885.4]
  wire  _T_1957; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293902.4]
  wire  _T_1958; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293903.4]
  wire  _T_1960; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293905.4]
  wire  _T_1962; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293907.4]
  wire [1:0] _T_1963; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293908.4]
  wire [1:0] _T_1964; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293909.4]
  wire  _T_1965; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293910.4]
  wire  _T_1966; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293912.4]
  wire  _T_1968; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293914.4]
  wire  _T_1970; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293916.4]
  wire  _T_1971; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293917.4]
  wire  _T_1972; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293922.4]
  wire  _T_1973; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293923.4]
  wire  _T_1974; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293924.4]
  wire  _T_1976; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293926.4]
  wire  _T_1977; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293927.4]
  wire  _T_1988; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293944.4]
  wire  _T_1989; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293945.4]
  wire  _T_1991; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293947.4]
  wire  _T_1993; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293949.4]
  wire [1:0] _T_1994; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293950.4]
  wire [1:0] _T_1995; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293951.4]
  wire  _T_1996; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293952.4]
  wire  _T_1997; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293954.4]
  wire  _T_1999; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293956.4]
  wire  _T_2001; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293958.4]
  wire  _T_2002; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293959.4]
  wire  _T_2003; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293964.4]
  wire  _T_2004; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293965.4]
  wire  _T_2005; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293966.4]
  wire  _T_2007; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293968.4]
  wire  _T_2008; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293969.4]
  wire  _T_2019; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293986.4]
  wire  _T_2020; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293987.4]
  wire  _T_2022; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293989.4]
  wire  _T_2024; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293991.4]
  wire [1:0] _T_2025; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293992.4]
  wire [1:0] _T_2026; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293993.4]
  wire  _T_2027; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293994.4]
  wire  _T_2028; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293996.4]
  wire  _T_2030; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293998.4]
  wire  _T_2032; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294000.4]
  wire  _T_2033; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294001.4]
  wire  _T_2034; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294006.4]
  wire  _T_2035; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294007.4]
  wire  _T_2036; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294008.4]
  wire  _T_2038; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294010.4]
  wire  _T_2039; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294011.4]
  wire  _T_2050; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294028.4]
  wire  _T_2051; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294029.4]
  wire  _T_2053; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294031.4]
  wire  _T_2055; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294033.4]
  wire [1:0] _T_2056; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294034.4]
  wire [1:0] _T_2057; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294035.4]
  wire  _T_2058; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294036.4]
  wire  _T_2059; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294038.4]
  wire  _T_2061; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294040.4]
  wire  _T_2063; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294042.4]
  wire  _T_2064; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294043.4]
  wire  _T_2065; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294048.4]
  wire  _T_2066; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294049.4]
  wire  _T_2067; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294050.4]
  wire  _T_2069; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294052.4]
  wire  _T_2070; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294053.4]
  wire  _T_2081; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294070.4]
  wire  _T_2082; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294071.4]
  wire  _T_2084; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294073.4]
  wire  _T_2086; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294075.4]
  wire [1:0] _T_2087; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294076.4]
  wire [1:0] _T_2088; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294077.4]
  wire  _T_2089; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294078.4]
  wire  _T_2090; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294080.4]
  wire  _T_2092; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294082.4]
  wire  _T_2094; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294084.4]
  wire  _T_2095; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294085.4]
  wire  _T_2096; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294090.4]
  wire  _T_2097; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294091.4]
  wire  _T_2098; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294092.4]
  wire  _T_2100; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294094.4]
  wire  _T_2101; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294095.4]
  wire  _T_2112; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294112.4]
  wire  _T_2113; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294113.4]
  wire  _T_2115; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294115.4]
  wire  _T_2117; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294117.4]
  wire [1:0] _T_2118; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294118.4]
  wire [1:0] _T_2119; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294119.4]
  wire  _T_2120; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294120.4]
  wire  _T_2121; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294122.4]
  wire  _T_2123; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294124.4]
  wire  _T_2125; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294126.4]
  wire  _T_2126; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294127.4]
  wire  _T_2127; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294132.4]
  wire  _T_2128; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294133.4]
  wire  _T_2129; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294134.4]
  wire  _T_2131; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294136.4]
  wire  _T_2132; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294137.4]
  wire  _T_2143; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294154.4]
  wire  _T_2144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294155.4]
  wire  _T_2146; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294157.4]
  wire  _T_2148; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294159.4]
  wire [1:0] _T_2149; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294160.4]
  wire [1:0] _T_2150; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294161.4]
  wire  _T_2151; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294162.4]
  wire  _T_2152; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294164.4]
  wire  _T_2154; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294166.4]
  wire  _T_2156; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294168.4]
  wire  _T_2157; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294169.4]
  wire  _T_2158; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294174.4]
  wire  _T_2159; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294175.4]
  wire  _T_2160; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294176.4]
  wire  _T_2162; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294178.4]
  wire  _T_2163; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294179.4]
  wire  _T_2174; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294196.4]
  wire  _T_2175; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294197.4]
  wire  _T_2177; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294199.4]
  wire  _T_2179; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294201.4]
  wire [1:0] _T_2180; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294202.4]
  wire [1:0] _T_2181; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294203.4]
  wire  _T_2182; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294204.4]
  wire  _T_2183; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294206.4]
  wire  _T_2185; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294208.4]
  wire  _T_2187; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294210.4]
  wire  _T_2188; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294211.4]
  wire  _T_2189; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294216.4]
  wire  _T_2190; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294217.4]
  wire  _T_2191; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294218.4]
  wire  _T_2193; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294220.4]
  wire  _T_2194; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294221.4]
  wire  _T_2205; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294238.4]
  wire  _T_2206; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294239.4]
  wire  _T_2208; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294241.4]
  wire  _T_2210; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294243.4]
  wire [1:0] _T_2211; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294244.4]
  wire [1:0] _T_2212; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294245.4]
  wire  _T_2213; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294246.4]
  wire  _T_2214; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294248.4]
  wire  _T_2216; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294250.4]
  wire  _T_2218; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294252.4]
  wire  _T_2219; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294253.4]
  wire  _T_2220; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294258.4]
  wire  _T_2221; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294259.4]
  wire  _T_2222; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294260.4]
  wire  _T_2224; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294262.4]
  wire  _T_2225; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294263.4]
  wire  _T_2236; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294280.4]
  wire  _T_2237; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294281.4]
  wire  _T_2239; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294283.4]
  wire  _T_2241; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294285.4]
  wire [1:0] _T_2242; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294286.4]
  wire [1:0] _T_2243; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294287.4]
  wire  _T_2244; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294288.4]
  wire  _T_2245; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294290.4]
  wire  _T_2247; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294292.4]
  wire  _T_2249; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294294.4]
  wire  _T_2250; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294295.4]
  wire  _T_2251; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294300.4]
  wire  _T_2252; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294301.4]
  wire  _T_2253; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294302.4]
  wire  _T_2255; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294304.4]
  wire  _T_2256; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294305.4]
  wire  _T_2267; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294322.4]
  wire  _T_2268; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294323.4]
  wire  _T_2270; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294325.4]
  wire  _T_2272; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294327.4]
  wire [1:0] _T_2273; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294328.4]
  wire [1:0] _T_2274; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294329.4]
  wire  _T_2275; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294330.4]
  wire  _T_2276; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294332.4]
  wire  _T_2278; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294334.4]
  wire  _T_2280; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294336.4]
  wire  _T_2281; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294337.4]
  wire  _T_2282; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294342.4]
  wire  _T_2283; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294343.4]
  wire  _T_2284; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294344.4]
  wire  _T_2286; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294346.4]
  wire  _T_2287; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294347.4]
  wire  _T_2298; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294364.4]
  wire  _T_2299; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294365.4]
  wire  _T_2301; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294367.4]
  wire  _T_2303; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294369.4]
  wire [1:0] _T_2304; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294370.4]
  wire [1:0] _T_2305; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294371.4]
  wire  _T_2306; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294372.4]
  wire  _T_2307; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294374.4]
  wire  _T_2309; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294376.4]
  wire  _T_2311; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294378.4]
  wire  _T_2312; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294379.4]
  wire  _T_2313; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294384.4]
  wire  _T_2314; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294385.4]
  wire  _T_2315; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294386.4]
  wire  _T_2317; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294388.4]
  wire  _T_2318; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294389.4]
  wire  _T_2329; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294406.4]
  wire  _T_2330; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294407.4]
  wire  _T_2332; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294409.4]
  wire  _T_2334; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294411.4]
  wire [1:0] _T_2335; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294412.4]
  wire [1:0] _T_2336; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294413.4]
  wire  _T_2337; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294414.4]
  wire  _T_2338; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294416.4]
  wire  _T_2340; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294418.4]
  wire  _T_2342; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294420.4]
  wire  _T_2343; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294421.4]
  wire  _T_2344; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294426.4]
  wire  _T_2345; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294427.4]
  wire  _T_2346; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294428.4]
  wire  _T_2348; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294430.4]
  wire  _T_2349; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294431.4]
  wire  _T_2360; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294448.4]
  wire  _T_2361; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294449.4]
  wire  _T_2363; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294451.4]
  wire  _T_2365; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294453.4]
  wire [1:0] _T_2366; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294454.4]
  wire [1:0] _T_2367; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294455.4]
  wire  _T_2368; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294456.4]
  wire  _T_2369; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294458.4]
  wire  _T_2371; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294460.4]
  wire  _T_2373; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294462.4]
  wire  _T_2374; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294463.4]
  wire  _T_2375; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294468.4]
  wire  _T_2376; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294469.4]
  wire  _T_2377; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294470.4]
  wire  _T_2379; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294472.4]
  wire  _T_2380; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294473.4]
  wire  _T_2391; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294490.4]
  wire  _T_2392; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294491.4]
  wire  _T_2394; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294493.4]
  wire  _T_2396; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294495.4]
  wire [1:0] _T_2397; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294496.4]
  wire [1:0] _T_2398; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294497.4]
  wire  _T_2399; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294498.4]
  wire  _T_2400; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294500.4]
  wire  _T_2402; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294502.4]
  wire  _T_2404; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294504.4]
  wire  _T_2405; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294505.4]
  wire  _T_2406; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294510.4]
  wire  _T_2407; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294511.4]
  wire  _T_2408; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294512.4]
  wire  _T_2410; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294514.4]
  wire  _T_2411; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294515.4]
  wire  _T_2422; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294532.4]
  wire  _T_2423; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294533.4]
  wire  _T_2425; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294535.4]
  wire  _T_2427; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294537.4]
  wire [1:0] _T_2428; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294538.4]
  wire [1:0] _T_2429; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294539.4]
  wire  _T_2430; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294540.4]
  wire  _T_2431; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294542.4]
  wire  _T_2433; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294544.4]
  wire  _T_2435; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294546.4]
  wire  _T_2436; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294547.4]
  wire  _T_2437; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294552.4]
  wire  _T_2438; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294553.4]
  wire  _T_2439; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294554.4]
  wire  _T_2441; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294556.4]
  wire  _T_2442; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294557.4]
  wire  _T_2453; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294574.4]
  wire  _T_2454; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294575.4]
  wire  _T_2456; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294577.4]
  wire  _T_2458; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294579.4]
  wire [1:0] _T_2459; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294580.4]
  wire [1:0] _T_2460; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294581.4]
  wire  _T_2461; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294582.4]
  wire  _T_2462; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294584.4]
  wire  _T_2464; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294586.4]
  wire  _T_2466; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294588.4]
  wire  _T_2467; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294589.4]
  wire  _T_2468; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294594.4]
  wire  _T_2469; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294595.4]
  wire  _T_2470; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294596.4]
  wire  _T_2472; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294598.4]
  wire  _T_2473; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294599.4]
  wire  _T_2484; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294616.4]
  wire  _T_2485; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294617.4]
  wire  _T_2487; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294619.4]
  wire  _T_2489; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294621.4]
  wire [1:0] _T_2490; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294622.4]
  wire [1:0] _T_2491; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294623.4]
  wire  _T_2492; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294624.4]
  wire  _T_2493; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294626.4]
  wire  _T_2495; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294628.4]
  wire  _T_2497; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294630.4]
  wire  _T_2498; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294631.4]
  wire  _T_2499; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294636.4]
  wire  _T_2500; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294637.4]
  wire  _T_2501; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294638.4]
  wire  _T_2503; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294640.4]
  wire  _T_2504; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294641.4]
  wire  _T_2515; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294658.4]
  wire  _T_2516; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294659.4]
  wire  _T_2518; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294661.4]
  wire  _T_2520; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294663.4]
  wire [1:0] _T_2521; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294664.4]
  wire [1:0] _T_2522; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294665.4]
  wire  _T_2523; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294666.4]
  wire  _T_2524; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294668.4]
  wire  _T_2526; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294670.4]
  wire  _T_2528; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294672.4]
  wire  _T_2529; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294673.4]
  wire  _T_2530; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294678.4]
  wire  _T_2531; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294679.4]
  wire  _T_2532; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294680.4]
  wire  _T_2534; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294682.4]
  wire  _T_2535; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294683.4]
  wire  _T_2546; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294700.4]
  wire  _T_2547; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294701.4]
  wire  _T_2549; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294703.4]
  wire  _T_2551; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294705.4]
  wire [1:0] _T_2552; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294706.4]
  wire [1:0] _T_2553; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294707.4]
  wire  _T_2554; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294708.4]
  wire  _T_2555; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294710.4]
  wire  _T_2557; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294712.4]
  wire  _T_2559; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294714.4]
  wire  _T_2560; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294715.4]
  wire  _T_2561; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294720.4]
  wire  _T_2562; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294721.4]
  wire  _T_2563; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294722.4]
  wire  _T_2565; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294724.4]
  wire  _T_2566; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294725.4]
  wire  _T_2577; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294742.4]
  wire  _T_2578; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294743.4]
  wire  _T_2580; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294745.4]
  wire  _T_2582; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294747.4]
  wire [1:0] _T_2583; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294748.4]
  wire [1:0] _T_2584; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294749.4]
  wire  _T_2585; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294750.4]
  wire  _T_2586; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294752.4]
  wire  _T_2588; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294754.4]
  wire  _T_2590; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294756.4]
  wire  _T_2591; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294757.4]
  wire  _T_2592; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294762.4]
  wire  _T_2593; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294763.4]
  wire  _T_2594; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294764.4]
  wire  _T_2596; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294766.4]
  wire  _T_2597; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294767.4]
  wire  _T_2608; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294784.4]
  wire  _T_2609; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294785.4]
  wire  _T_2611; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294787.4]
  wire  _T_2613; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294789.4]
  wire [1:0] _T_2614; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294790.4]
  wire [1:0] _T_2615; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294791.4]
  wire  _T_2616; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294792.4]
  wire  _T_2617; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294794.4]
  wire  _T_2619; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294796.4]
  wire  _T_2621; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294798.4]
  wire  _T_2622; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294799.4]
  wire  _T_2623; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294804.4]
  wire  _T_2624; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294805.4]
  wire  _T_2625; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294806.4]
  wire  _T_2627; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294808.4]
  wire  _T_2628; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294809.4]
  wire  _T_2639; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294826.4]
  wire  _T_2640; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294827.4]
  wire  _T_2642; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294829.4]
  wire  _T_2644; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294831.4]
  wire [1:0] _T_2645; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294832.4]
  wire [1:0] _T_2646; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294833.4]
  wire  _T_2647; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294834.4]
  wire  _T_2648; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294836.4]
  wire  _T_2650; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294838.4]
  wire  _T_2652; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294840.4]
  wire  _T_2653; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294841.4]
  wire  _T_2654; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294846.4]
  wire  _T_2655; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294847.4]
  wire  _T_2656; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294848.4]
  wire  _T_2658; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294850.4]
  wire  _T_2659; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294851.4]
  wire  _T_2670; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294868.4]
  wire  _T_2671; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294869.4]
  wire  _T_2673; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294871.4]
  wire  _T_2675; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294873.4]
  wire [1:0] _T_2676; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294874.4]
  wire [1:0] _T_2677; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294875.4]
  wire  _T_2678; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294876.4]
  wire  _T_2679; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294878.4]
  wire  _T_2681; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294880.4]
  wire  _T_2683; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294882.4]
  wire  _T_2684; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294883.4]
  wire  _T_2685; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294888.4]
  wire  _T_2686; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294889.4]
  wire  _T_2687; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294890.4]
  wire  _T_2689; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294892.4]
  wire  _T_2690; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294893.4]
  wire  _T_2701; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294910.4]
  wire  _T_2702; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294911.4]
  wire  _T_2704; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294913.4]
  wire  _T_2706; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294915.4]
  wire [1:0] _T_2707; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294916.4]
  wire [1:0] _T_2708; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294917.4]
  wire  _T_2709; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294918.4]
  wire  _T_2710; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294920.4]
  wire  _T_2712; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294922.4]
  wire  _T_2714; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294924.4]
  wire  _T_2715; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294925.4]
  wire  _T_2716; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294930.4]
  wire  _T_2717; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294931.4]
  wire  _T_2718; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294932.4]
  wire  _T_2720; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294934.4]
  wire  _T_2721; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294935.4]
  wire  _T_2732; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294952.4]
  wire  _T_2733; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294953.4]
  wire  _T_2735; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294955.4]
  wire  _T_2737; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294957.4]
  wire [1:0] _T_2738; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294958.4]
  wire [1:0] _T_2739; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294959.4]
  wire  _T_2740; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294960.4]
  wire  _T_2741; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294962.4]
  wire  _T_2743; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294964.4]
  wire  _T_2745; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294966.4]
  wire  _T_2746; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294967.4]
  wire  _T_2747; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294972.4]
  wire  _T_2748; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294973.4]
  wire  _T_2749; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294974.4]
  wire  _T_2751; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294976.4]
  wire  _T_2752; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294977.4]
  wire  _T_2763; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294994.4]
  wire  _T_2764; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294995.4]
  wire  _T_2766; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294997.4]
  wire  _T_2768; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294999.4]
  wire [1:0] _T_2769; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295000.4]
  wire [1:0] _T_2770; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295001.4]
  wire  _T_2771; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295002.4]
  wire  _T_2772; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295004.4]
  wire  _T_2774; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295006.4]
  wire  _T_2776; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295008.4]
  wire  _T_2777; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295009.4]
  wire  _T_2778; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295014.4]
  wire  _T_2779; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295015.4]
  wire  _T_2780; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295016.4]
  wire  _T_2782; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295018.4]
  wire  _T_2783; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295019.4]
  wire  _T_2794; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295036.4]
  wire  _T_2795; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295037.4]
  wire  _T_2797; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295039.4]
  wire  _T_2799; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295041.4]
  wire [1:0] _T_2800; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295042.4]
  wire [1:0] _T_2801; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295043.4]
  wire  _T_2802; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295044.4]
  wire  _T_2803; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295046.4]
  wire  _T_2805; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295048.4]
  wire  _T_2807; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295050.4]
  wire  _T_2808; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295051.4]
  wire  _T_2809; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295056.4]
  wire  _T_2810; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295057.4]
  wire  _T_2811; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295058.4]
  wire  _T_2813; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295060.4]
  wire  _T_2814; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295061.4]
  wire  _T_2825; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295078.4]
  wire  _T_2826; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295079.4]
  wire  _T_2828; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295081.4]
  wire  _T_2830; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295083.4]
  wire [1:0] _T_2831; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295084.4]
  wire [1:0] _T_2832; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295085.4]
  wire  _T_2833; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295086.4]
  wire  _T_2834; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295088.4]
  wire  _T_2836; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295090.4]
  wire  _T_2838; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295092.4]
  wire  _T_2839; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295093.4]
  wire  _T_2840; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295098.4]
  wire  _T_2841; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295099.4]
  wire  _T_2842; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295100.4]
  wire  _T_2844; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295102.4]
  wire  _T_2845; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295103.4]
  wire  _T_2856; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295120.4]
  wire  _T_2857; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295121.4]
  wire  _T_2859; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295123.4]
  wire  _T_2861; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295125.4]
  wire [1:0] _T_2862; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295126.4]
  wire [1:0] _T_2863; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295127.4]
  wire  _T_2864; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295128.4]
  wire  _T_2865; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295130.4]
  wire  _T_2867; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295132.4]
  wire  _T_2869; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295134.4]
  wire  _T_2870; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295135.4]
  wire  _T_2871; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295140.4]
  wire  _T_2872; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295141.4]
  wire  _T_2873; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295142.4]
  wire  _T_2875; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295144.4]
  wire  _T_2876; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295145.4]
  wire  _T_2887; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295162.4]
  wire  _T_2888; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295163.4]
  wire  _T_2890; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295165.4]
  wire  _T_2892; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295167.4]
  wire [1:0] _T_2893; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295168.4]
  wire [1:0] _T_2894; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295169.4]
  wire  _T_2895; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295170.4]
  wire  _T_2896; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295172.4]
  wire  _T_2898; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295174.4]
  wire  _T_2900; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295176.4]
  wire  _T_2901; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295177.4]
  wire  _T_2902; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295182.4]
  wire  _T_2903; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295183.4]
  wire  _T_2904; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295184.4]
  wire  _T_2906; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295186.4]
  wire  _T_2907; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295187.4]
  wire  _T_2918; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295204.4]
  wire  _T_2919; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295205.4]
  wire  _T_2921; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295207.4]
  wire  _T_2923; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295209.4]
  wire [1:0] _T_2924; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295210.4]
  wire [1:0] _T_2925; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295211.4]
  wire  _T_2926; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295212.4]
  wire  _T_2927; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295214.4]
  wire  _T_2929; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295216.4]
  wire  _T_2931; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295218.4]
  wire  _T_2932; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295219.4]
  wire  _T_2933; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295224.4]
  wire  _T_2934; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295225.4]
  wire  _T_2935; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295226.4]
  wire  _T_2937; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295228.4]
  wire  _T_2938; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295229.4]
  wire  _T_2949; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295246.4]
  wire  _T_2950; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295247.4]
  wire  _T_2952; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295249.4]
  wire  _T_2954; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295251.4]
  wire [1:0] _T_2955; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295252.4]
  wire [1:0] _T_2956; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295253.4]
  wire  _T_2957; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295254.4]
  wire  _T_2958; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295256.4]
  wire  _T_2960; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295258.4]
  wire  _T_2962; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295260.4]
  wire  _T_2963; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295261.4]
  wire  _T_2964; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295266.4]
  wire  _T_2965; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295267.4]
  wire  _T_2966; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295268.4]
  wire  _T_2968; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295270.4]
  wire  _T_2969; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295271.4]
  wire  _T_2980; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295288.4]
  wire  _T_2981; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295289.4]
  wire  _T_2983; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295291.4]
  wire  _T_2985; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295293.4]
  wire [1:0] _T_2986; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295294.4]
  wire [1:0] _T_2987; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295295.4]
  wire  _T_2988; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295296.4]
  wire  _T_2989; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295298.4]
  wire  _T_2991; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295300.4]
  wire  _T_2993; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295302.4]
  wire  _T_2994; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295303.4]
  wire  _T_2995; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295308.4]
  wire  _T_2996; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295309.4]
  wire  _T_2997; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295310.4]
  wire  _T_2999; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295312.4]
  wire  _T_3000; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295313.4]
  wire  _T_3011; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295330.4]
  wire  _T_3012; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295331.4]
  wire  _T_3014; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295333.4]
  wire  _T_3016; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295335.4]
  wire [1:0] _T_3017; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295336.4]
  wire [1:0] _T_3018; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295337.4]
  wire  _T_3019; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295338.4]
  wire  _T_3020; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295340.4]
  wire  _T_3022; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295342.4]
  wire  _T_3024; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295344.4]
  wire  _T_3025; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295345.4]
  wire  _T_3026; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295350.4]
  wire  _T_3027; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295351.4]
  wire  _T_3028; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295352.4]
  wire  _T_3030; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295354.4]
  wire  _T_3031; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295355.4]
  wire  _T_3042; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295372.4]
  wire  _T_3043; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295373.4]
  wire  _T_3045; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295375.4]
  wire  _T_3047; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295377.4]
  wire [1:0] _T_3048; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295378.4]
  wire [1:0] _T_3049; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295379.4]
  wire  _T_3050; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295380.4]
  wire  _T_3051; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295382.4]
  wire  _T_3053; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295384.4]
  wire  _T_3055; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295386.4]
  wire  _T_3056; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295387.4]
  wire  _T_3057; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295392.4]
  wire  _T_3058; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295393.4]
  wire  _T_3059; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295394.4]
  wire  _T_3061; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295396.4]
  wire  _T_3062; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295397.4]
  wire  _T_3073; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295414.4]
  wire  _T_3074; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295415.4]
  wire  _T_3076; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295417.4]
  wire  _T_3078; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295419.4]
  wire [1:0] _T_3079; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295420.4]
  wire [1:0] _T_3080; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295421.4]
  wire  _T_3081; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295422.4]
  wire  _T_3082; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295424.4]
  wire  _T_3084; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295426.4]
  wire  _T_3086; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295428.4]
  wire  _T_3087; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295429.4]
  wire  _T_3088; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295434.4]
  wire  _T_3089; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295435.4]
  wire  _T_3090; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295436.4]
  wire  _T_3092; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295438.4]
  wire  _T_3093; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295439.4]
  wire  _T_3104; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295456.4]
  wire  _T_3105; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295457.4]
  wire  _T_3107; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295459.4]
  wire  _T_3109; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295461.4]
  wire [1:0] _T_3110; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295462.4]
  wire [1:0] _T_3111; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295463.4]
  wire  _T_3112; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295464.4]
  wire  _T_3113; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295466.4]
  wire  _T_3115; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295468.4]
  wire  _T_3117; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295470.4]
  wire  _T_3118; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295471.4]
  wire  _T_3119; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295476.4]
  wire  _T_3120; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295477.4]
  wire  _T_3121; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295478.4]
  wire  _T_3123; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295480.4]
  wire  _T_3124; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295481.4]
  Queue_44 Queue ( // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292519.4]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_strb(Queue_io_enq_bits_strb),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_strb(Queue_io_deq_bits_strb),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_45 Queue_1 ( // @[Decoupled.scala 293:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292534.4]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_wen(Queue_1_io_enq_bits_wen),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_1_io_deq_bits_qos),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_wen(Queue_1_io_deq_bits_wen)
  );
  assign _T_887 = auto_in_a_bits_opcode[2]; // @[Edges.scala 92:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292466.4]
  assign _T_888 = _T_887 == 1'h0; // @[Edges.scala 92:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292467.4]
  assign _GEN_132 = 7'h2 == auto_in_a_bits_source ? _T_1177 : _T_1146; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_133 = 7'h3 == auto_in_a_bits_source ? _T_1177 : _GEN_132; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_134 = 7'h4 == auto_in_a_bits_source ? _T_1208 : _GEN_133; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_135 = 7'h5 == auto_in_a_bits_source ? _T_1208 : _GEN_134; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_136 = 7'h6 == auto_in_a_bits_source ? _T_1239 : _GEN_135; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_137 = 7'h7 == auto_in_a_bits_source ? _T_1239 : _GEN_136; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_138 = 7'h8 == auto_in_a_bits_source ? _T_1270 : _GEN_137; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_139 = 7'h9 == auto_in_a_bits_source ? _T_1270 : _GEN_138; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_140 = 7'ha == auto_in_a_bits_source ? _T_1301 : _GEN_139; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_141 = 7'hb == auto_in_a_bits_source ? _T_1301 : _GEN_140; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_142 = 7'hc == auto_in_a_bits_source ? _T_1332 : _GEN_141; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_143 = 7'hd == auto_in_a_bits_source ? _T_1332 : _GEN_142; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_144 = 7'he == auto_in_a_bits_source ? _T_1363 : _GEN_143; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_145 = 7'hf == auto_in_a_bits_source ? _T_1363 : _GEN_144; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_146 = 7'h10 == auto_in_a_bits_source ? _T_1394 : _GEN_145; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_147 = 7'h11 == auto_in_a_bits_source ? _T_1394 : _GEN_146; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_148 = 7'h12 == auto_in_a_bits_source ? _T_1425 : _GEN_147; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_149 = 7'h13 == auto_in_a_bits_source ? _T_1425 : _GEN_148; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_150 = 7'h14 == auto_in_a_bits_source ? _T_1456 : _GEN_149; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_151 = 7'h15 == auto_in_a_bits_source ? _T_1456 : _GEN_150; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_152 = 7'h16 == auto_in_a_bits_source ? _T_1487 : _GEN_151; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_153 = 7'h17 == auto_in_a_bits_source ? _T_1487 : _GEN_152; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_154 = 7'h18 == auto_in_a_bits_source ? _T_1518 : _GEN_153; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_155 = 7'h19 == auto_in_a_bits_source ? _T_1518 : _GEN_154; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_156 = 7'h1a == auto_in_a_bits_source ? _T_1549 : _GEN_155; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_157 = 7'h1b == auto_in_a_bits_source ? _T_1549 : _GEN_156; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_158 = 7'h1c == auto_in_a_bits_source ? _T_1580 : _GEN_157; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_159 = 7'h1d == auto_in_a_bits_source ? _T_1580 : _GEN_158; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_160 = 7'h1e == auto_in_a_bits_source ? _T_1611 : _GEN_159; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_161 = 7'h1f == auto_in_a_bits_source ? _T_1611 : _GEN_160; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_162 = 7'h20 == auto_in_a_bits_source ? _T_1642 : _GEN_161; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_163 = 7'h21 == auto_in_a_bits_source ? _T_1642 : _GEN_162; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_164 = 7'h22 == auto_in_a_bits_source ? _T_1673 : _GEN_163; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_165 = 7'h23 == auto_in_a_bits_source ? _T_1673 : _GEN_164; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_166 = 7'h24 == auto_in_a_bits_source ? _T_1704 : _GEN_165; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_167 = 7'h25 == auto_in_a_bits_source ? _T_1704 : _GEN_166; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_168 = 7'h26 == auto_in_a_bits_source ? _T_1735 : _GEN_167; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_169 = 7'h27 == auto_in_a_bits_source ? _T_1735 : _GEN_168; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_170 = 7'h28 == auto_in_a_bits_source ? _T_1766 : _GEN_169; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_171 = 7'h29 == auto_in_a_bits_source ? _T_1766 : _GEN_170; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_172 = 7'h2a == auto_in_a_bits_source ? _T_1797 : _GEN_171; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_173 = 7'h2b == auto_in_a_bits_source ? _T_1797 : _GEN_172; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_174 = 7'h2c == auto_in_a_bits_source ? _T_1828 : _GEN_173; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_175 = 7'h2d == auto_in_a_bits_source ? _T_1828 : _GEN_174; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_176 = 7'h2e == auto_in_a_bits_source ? _T_1859 : _GEN_175; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_177 = 7'h2f == auto_in_a_bits_source ? _T_1859 : _GEN_176; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_178 = 7'h30 == auto_in_a_bits_source ? _T_1890 : _GEN_177; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_179 = 7'h31 == auto_in_a_bits_source ? _T_1890 : _GEN_178; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_180 = 7'h32 == auto_in_a_bits_source ? _T_1921 : _GEN_179; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_181 = 7'h33 == auto_in_a_bits_source ? _T_1921 : _GEN_180; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_182 = 7'h34 == auto_in_a_bits_source ? _T_1952 : _GEN_181; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_183 = 7'h35 == auto_in_a_bits_source ? _T_1952 : _GEN_182; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_184 = 7'h36 == auto_in_a_bits_source ? _T_1983 : _GEN_183; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_185 = 7'h37 == auto_in_a_bits_source ? _T_1983 : _GEN_184; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_186 = 7'h38 == auto_in_a_bits_source ? _T_2014 : _GEN_185; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_187 = 7'h39 == auto_in_a_bits_source ? _T_2014 : _GEN_186; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_188 = 7'h3a == auto_in_a_bits_source ? _T_2045 : _GEN_187; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_189 = 7'h3b == auto_in_a_bits_source ? _T_2045 : _GEN_188; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_190 = 7'h3c == auto_in_a_bits_source ? _T_2076 : _GEN_189; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_191 = 7'h3d == auto_in_a_bits_source ? _T_2076 : _GEN_190; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_192 = 7'h3e == auto_in_a_bits_source ? _T_2107 : _GEN_191; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_193 = 7'h3f == auto_in_a_bits_source ? _T_2107 : _GEN_192; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_194 = 7'h40 == auto_in_a_bits_source ? _T_2138 : _GEN_193; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_195 = 7'h41 == auto_in_a_bits_source ? _T_2138 : _GEN_194; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_196 = 7'h42 == auto_in_a_bits_source ? _T_2169 : _GEN_195; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_197 = 7'h43 == auto_in_a_bits_source ? _T_2169 : _GEN_196; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_198 = 7'h44 == auto_in_a_bits_source ? _T_2200 : _GEN_197; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_199 = 7'h45 == auto_in_a_bits_source ? _T_2200 : _GEN_198; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_200 = 7'h46 == auto_in_a_bits_source ? _T_2231 : _GEN_199; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_201 = 7'h47 == auto_in_a_bits_source ? _T_2231 : _GEN_200; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_202 = 7'h48 == auto_in_a_bits_source ? _T_2262 : _GEN_201; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_203 = 7'h49 == auto_in_a_bits_source ? _T_2262 : _GEN_202; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_204 = 7'h4a == auto_in_a_bits_source ? _T_2293 : _GEN_203; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_205 = 7'h4b == auto_in_a_bits_source ? _T_2293 : _GEN_204; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_206 = 7'h4c == auto_in_a_bits_source ? _T_2324 : _GEN_205; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_207 = 7'h4d == auto_in_a_bits_source ? _T_2324 : _GEN_206; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_208 = 7'h4e == auto_in_a_bits_source ? _T_2355 : _GEN_207; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_209 = 7'h4f == auto_in_a_bits_source ? _T_2355 : _GEN_208; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_210 = 7'h50 == auto_in_a_bits_source ? _T_2386 : _GEN_209; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_211 = 7'h51 == auto_in_a_bits_source ? _T_2386 : _GEN_210; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_212 = 7'h52 == auto_in_a_bits_source ? _T_2417 : _GEN_211; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_213 = 7'h53 == auto_in_a_bits_source ? _T_2417 : _GEN_212; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_214 = 7'h54 == auto_in_a_bits_source ? _T_2448 : _GEN_213; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_215 = 7'h55 == auto_in_a_bits_source ? _T_2448 : _GEN_214; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_216 = 7'h56 == auto_in_a_bits_source ? _T_2479 : _GEN_215; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_217 = 7'h57 == auto_in_a_bits_source ? _T_2479 : _GEN_216; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_218 = 7'h58 == auto_in_a_bits_source ? _T_2510 : _GEN_217; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_219 = 7'h59 == auto_in_a_bits_source ? _T_2510 : _GEN_218; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_220 = 7'h5a == auto_in_a_bits_source ? _T_2541 : _GEN_219; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_221 = 7'h5b == auto_in_a_bits_source ? _T_2541 : _GEN_220; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_222 = 7'h5c == auto_in_a_bits_source ? _T_2572 : _GEN_221; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_223 = 7'h5d == auto_in_a_bits_source ? _T_2572 : _GEN_222; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_224 = 7'h5e == auto_in_a_bits_source ? _T_2603 : _GEN_223; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_225 = 7'h5f == auto_in_a_bits_source ? _T_2603 : _GEN_224; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_226 = 7'h60 == auto_in_a_bits_source ? _T_2634 : _GEN_225; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_227 = 7'h61 == auto_in_a_bits_source ? _T_2634 : _GEN_226; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_228 = 7'h62 == auto_in_a_bits_source ? _T_2665 : _GEN_227; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_229 = 7'h63 == auto_in_a_bits_source ? _T_2665 : _GEN_228; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_230 = 7'h64 == auto_in_a_bits_source ? _T_2696 : _GEN_229; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_231 = 7'h65 == auto_in_a_bits_source ? _T_2696 : _GEN_230; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_232 = 7'h66 == auto_in_a_bits_source ? _T_2727 : _GEN_231; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_233 = 7'h67 == auto_in_a_bits_source ? _T_2727 : _GEN_232; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_234 = 7'h68 == auto_in_a_bits_source ? _T_2758 : _GEN_233; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_235 = 7'h69 == auto_in_a_bits_source ? _T_2758 : _GEN_234; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_236 = 7'h6a == auto_in_a_bits_source ? _T_2789 : _GEN_235; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_237 = 7'h6b == auto_in_a_bits_source ? _T_2789 : _GEN_236; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_238 = 7'h6c == auto_in_a_bits_source ? _T_2820 : _GEN_237; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_239 = 7'h6d == auto_in_a_bits_source ? _T_2820 : _GEN_238; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_240 = 7'h6e == auto_in_a_bits_source ? _T_2851 : _GEN_239; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_241 = 7'h6f == auto_in_a_bits_source ? _T_2851 : _GEN_240; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_242 = 7'h70 == auto_in_a_bits_source ? _T_2882 : _GEN_241; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_243 = 7'h71 == auto_in_a_bits_source ? _T_2882 : _GEN_242; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_244 = 7'h72 == auto_in_a_bits_source ? _T_2913 : _GEN_243; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_245 = 7'h73 == auto_in_a_bits_source ? _T_2913 : _GEN_244; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_246 = 7'h74 == auto_in_a_bits_source ? _T_2944 : _GEN_245; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_247 = 7'h75 == auto_in_a_bits_source ? _T_2944 : _GEN_246; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_248 = 7'h76 == auto_in_a_bits_source ? _T_2975 : _GEN_247; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_249 = 7'h77 == auto_in_a_bits_source ? _T_2975 : _GEN_248; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_250 = 7'h78 == auto_in_a_bits_source ? _T_3006 : _GEN_249; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_251 = 7'h79 == auto_in_a_bits_source ? _T_3006 : _GEN_250; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_252 = 7'h7a == auto_in_a_bits_source ? _T_3037 : _GEN_251; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_253 = 7'h7b == auto_in_a_bits_source ? _T_3037 : _GEN_252; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_254 = 7'h7c == auto_in_a_bits_source ? _T_3068 : _GEN_253; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_255 = 7'h7d == auto_in_a_bits_source ? _T_3068 : _GEN_254; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_256 = 7'h7e == auto_in_a_bits_source ? _T_3099 : _GEN_255; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _GEN_257 = 7'h7f == auto_in_a_bits_source ? _T_3099 : _GEN_256; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _T_903 = _T_899 == 4'h0; // @[Edges.scala 231:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292481.4]
  assign _T_969 = _GEN_257 & _T_903; // @[ToAXI4.scala 176:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292597.4]
  assign _T_970 = _T_969 == 1'h0; // @[ToAXI4.scala 177:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292598.4]
  assign _T_930_ready = Queue_1_io_enq_ready; // @[ToAXI4.scala 146:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292515.4 Decoupled.scala 296:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292549.4]
  assign _T_971 = _T_957 | _T_930_ready; // @[ToAXI4.scala 177:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292599.4]
  assign _T_933_ready = Queue_io_enq_ready; // @[ToAXI4.scala 147:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292517.4 Decoupled.scala 296:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292526.4]
  assign _T_972 = _T_971 & _T_933_ready; // @[ToAXI4.scala 177:70:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292600.4]
  assign _T_973 = _T_888 ? _T_972 : _T_930_ready; // @[ToAXI4.scala 177:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292601.4]
  assign _T_974 = _T_970 & _T_973; // @[ToAXI4.scala 177:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292602.4]
  assign _T_889 = _T_974 & auto_in_a_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292468.4]
  assign _T_891 = 14'h7f << auto_in_a_bits_size; // @[package.scala 185:77:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292470.4]
  assign _T_892 = _T_891[6:0]; // @[package.scala 185:82:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292471.4]
  assign _T_893 = ~ _T_892; // @[package.scala 185:46:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292472.4]
  assign _T_894 = _T_893[6:3]; // @[Edges.scala 220:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292473.4]
  assign _T_897 = _T_888 ? _T_894 : 4'h0; // @[Edges.scala 221:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292476.4]
  assign _T_900 = _T_899 - 4'h1; // @[Edges.scala 230:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292478.4]
  assign _T_901 = $unsigned(_T_900); // @[Edges.scala 230:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292479.4]
  assign _T_902 = _T_901[3:0]; // @[Edges.scala 230:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292480.4]
  assign _T_904 = _T_899 == 4'h1; // @[Edges.scala 232:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292482.4]
  assign _T_905 = _T_897 == 4'h0; // @[Edges.scala 232:47:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292483.4]
  assign _T_906 = _T_904 | _T_905; // @[Edges.scala 232:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292484.4]
  assign _GEN_325 = {{7'd0}, auto_in_a_bits_size}; // @[ToAXI4.scala 134:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292509.4]
  assign _T_920 = _GEN_325 << 7; // @[ToAXI4.scala 134:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292509.4]
  assign _GEN_326 = {{3'd0}, auto_in_a_bits_source}; // @[ToAXI4.scala 134:45:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292510.4]
  assign _T_921 = _GEN_326 | _T_920; // @[ToAXI4.scala 134:45:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292510.4]
  assign _T_922 = auto_out_r_bits_user[6:0]; // @[ToAXI4.scala 137:50:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292511.4]
  assign _T_923 = auto_out_r_bits_user[9:7]; // @[ToAXI4.scala 138:50:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292512.4]
  assign _T_924 = auto_out_b_bits_user[6:0]; // @[ToAXI4.scala 141:50:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292513.4]
  assign _T_925 = auto_out_b_bits_user[9:7]; // @[ToAXI4.scala 142:50:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292514.4]
  assign _T_948_bits_wen = Queue_1_io_deq_bits_wen; // @[Decoupled.scala 314:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292550.4 Decoupled.scala 315:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292551.4]
  assign _T_952 = _T_948_bits_wen == 1'h0; // @[ToAXI4.scala 154:42:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292566.4]
  assign _T_948_valid = Queue_1_io_deq_valid; // @[Decoupled.scala 314:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292550.4 Decoupled.scala 316:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292562.4]
  assign _T_959 = _T_906 == 1'h0; // @[ToAXI4.scala 161:38:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292576.6]
  assign _GEN_4 = 7'h2 == auto_in_a_bits_source ? 6'h1 : 6'h0; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_5 = 7'h3 == auto_in_a_bits_source ? 6'h1 : _GEN_4; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_6 = 7'h4 == auto_in_a_bits_source ? 6'h2 : _GEN_5; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_7 = 7'h5 == auto_in_a_bits_source ? 6'h2 : _GEN_6; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_8 = 7'h6 == auto_in_a_bits_source ? 6'h3 : _GEN_7; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_9 = 7'h7 == auto_in_a_bits_source ? 6'h3 : _GEN_8; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_10 = 7'h8 == auto_in_a_bits_source ? 6'h4 : _GEN_9; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_11 = 7'h9 == auto_in_a_bits_source ? 6'h4 : _GEN_10; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_12 = 7'ha == auto_in_a_bits_source ? 6'h5 : _GEN_11; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_13 = 7'hb == auto_in_a_bits_source ? 6'h5 : _GEN_12; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_14 = 7'hc == auto_in_a_bits_source ? 6'h6 : _GEN_13; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_15 = 7'hd == auto_in_a_bits_source ? 6'h6 : _GEN_14; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_16 = 7'he == auto_in_a_bits_source ? 6'h7 : _GEN_15; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_17 = 7'hf == auto_in_a_bits_source ? 6'h7 : _GEN_16; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_18 = 7'h10 == auto_in_a_bits_source ? 6'h8 : _GEN_17; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_19 = 7'h11 == auto_in_a_bits_source ? 6'h8 : _GEN_18; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_20 = 7'h12 == auto_in_a_bits_source ? 6'h9 : _GEN_19; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_21 = 7'h13 == auto_in_a_bits_source ? 6'h9 : _GEN_20; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_22 = 7'h14 == auto_in_a_bits_source ? 6'ha : _GEN_21; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_23 = 7'h15 == auto_in_a_bits_source ? 6'ha : _GEN_22; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_24 = 7'h16 == auto_in_a_bits_source ? 6'hb : _GEN_23; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_25 = 7'h17 == auto_in_a_bits_source ? 6'hb : _GEN_24; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_26 = 7'h18 == auto_in_a_bits_source ? 6'hc : _GEN_25; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_27 = 7'h19 == auto_in_a_bits_source ? 6'hc : _GEN_26; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_28 = 7'h1a == auto_in_a_bits_source ? 6'hd : _GEN_27; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_29 = 7'h1b == auto_in_a_bits_source ? 6'hd : _GEN_28; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_30 = 7'h1c == auto_in_a_bits_source ? 6'he : _GEN_29; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_31 = 7'h1d == auto_in_a_bits_source ? 6'he : _GEN_30; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_32 = 7'h1e == auto_in_a_bits_source ? 6'hf : _GEN_31; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_33 = 7'h1f == auto_in_a_bits_source ? 6'hf : _GEN_32; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_34 = 7'h20 == auto_in_a_bits_source ? 6'h10 : _GEN_33; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_35 = 7'h21 == auto_in_a_bits_source ? 6'h10 : _GEN_34; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_36 = 7'h22 == auto_in_a_bits_source ? 6'h11 : _GEN_35; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_37 = 7'h23 == auto_in_a_bits_source ? 6'h11 : _GEN_36; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_38 = 7'h24 == auto_in_a_bits_source ? 6'h12 : _GEN_37; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_39 = 7'h25 == auto_in_a_bits_source ? 6'h12 : _GEN_38; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_40 = 7'h26 == auto_in_a_bits_source ? 6'h13 : _GEN_39; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_41 = 7'h27 == auto_in_a_bits_source ? 6'h13 : _GEN_40; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_42 = 7'h28 == auto_in_a_bits_source ? 6'h14 : _GEN_41; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_43 = 7'h29 == auto_in_a_bits_source ? 6'h14 : _GEN_42; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_44 = 7'h2a == auto_in_a_bits_source ? 6'h15 : _GEN_43; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_45 = 7'h2b == auto_in_a_bits_source ? 6'h15 : _GEN_44; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_46 = 7'h2c == auto_in_a_bits_source ? 6'h16 : _GEN_45; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_47 = 7'h2d == auto_in_a_bits_source ? 6'h16 : _GEN_46; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_48 = 7'h2e == auto_in_a_bits_source ? 6'h17 : _GEN_47; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_49 = 7'h2f == auto_in_a_bits_source ? 6'h17 : _GEN_48; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_50 = 7'h30 == auto_in_a_bits_source ? 6'h18 : _GEN_49; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_51 = 7'h31 == auto_in_a_bits_source ? 6'h18 : _GEN_50; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_52 = 7'h32 == auto_in_a_bits_source ? 6'h19 : _GEN_51; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_53 = 7'h33 == auto_in_a_bits_source ? 6'h19 : _GEN_52; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_54 = 7'h34 == auto_in_a_bits_source ? 6'h1a : _GEN_53; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_55 = 7'h35 == auto_in_a_bits_source ? 6'h1a : _GEN_54; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_56 = 7'h36 == auto_in_a_bits_source ? 6'h1b : _GEN_55; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_57 = 7'h37 == auto_in_a_bits_source ? 6'h1b : _GEN_56; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_58 = 7'h38 == auto_in_a_bits_source ? 6'h1c : _GEN_57; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_59 = 7'h39 == auto_in_a_bits_source ? 6'h1c : _GEN_58; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_60 = 7'h3a == auto_in_a_bits_source ? 6'h1d : _GEN_59; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_61 = 7'h3b == auto_in_a_bits_source ? 6'h1d : _GEN_60; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_62 = 7'h3c == auto_in_a_bits_source ? 6'h1e : _GEN_61; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_63 = 7'h3d == auto_in_a_bits_source ? 6'h1e : _GEN_62; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_64 = 7'h3e == auto_in_a_bits_source ? 6'h1f : _GEN_63; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_65 = 7'h3f == auto_in_a_bits_source ? 6'h1f : _GEN_64; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_66 = 7'h40 == auto_in_a_bits_source ? 6'h20 : _GEN_65; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_67 = 7'h41 == auto_in_a_bits_source ? 6'h20 : _GEN_66; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_68 = 7'h42 == auto_in_a_bits_source ? 6'h21 : _GEN_67; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_69 = 7'h43 == auto_in_a_bits_source ? 6'h21 : _GEN_68; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_70 = 7'h44 == auto_in_a_bits_source ? 6'h22 : _GEN_69; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_71 = 7'h45 == auto_in_a_bits_source ? 6'h22 : _GEN_70; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_72 = 7'h46 == auto_in_a_bits_source ? 6'h23 : _GEN_71; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_73 = 7'h47 == auto_in_a_bits_source ? 6'h23 : _GEN_72; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_74 = 7'h48 == auto_in_a_bits_source ? 6'h24 : _GEN_73; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_75 = 7'h49 == auto_in_a_bits_source ? 6'h24 : _GEN_74; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_76 = 7'h4a == auto_in_a_bits_source ? 6'h25 : _GEN_75; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_77 = 7'h4b == auto_in_a_bits_source ? 6'h25 : _GEN_76; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_78 = 7'h4c == auto_in_a_bits_source ? 6'h26 : _GEN_77; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_79 = 7'h4d == auto_in_a_bits_source ? 6'h26 : _GEN_78; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_80 = 7'h4e == auto_in_a_bits_source ? 6'h27 : _GEN_79; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_81 = 7'h4f == auto_in_a_bits_source ? 6'h27 : _GEN_80; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_82 = 7'h50 == auto_in_a_bits_source ? 6'h28 : _GEN_81; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_83 = 7'h51 == auto_in_a_bits_source ? 6'h28 : _GEN_82; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_84 = 7'h52 == auto_in_a_bits_source ? 6'h29 : _GEN_83; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_85 = 7'h53 == auto_in_a_bits_source ? 6'h29 : _GEN_84; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_86 = 7'h54 == auto_in_a_bits_source ? 6'h2a : _GEN_85; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_87 = 7'h55 == auto_in_a_bits_source ? 6'h2a : _GEN_86; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_88 = 7'h56 == auto_in_a_bits_source ? 6'h2b : _GEN_87; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_89 = 7'h57 == auto_in_a_bits_source ? 6'h2b : _GEN_88; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_90 = 7'h58 == auto_in_a_bits_source ? 6'h2c : _GEN_89; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_91 = 7'h59 == auto_in_a_bits_source ? 6'h2c : _GEN_90; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_92 = 7'h5a == auto_in_a_bits_source ? 6'h2d : _GEN_91; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_93 = 7'h5b == auto_in_a_bits_source ? 6'h2d : _GEN_92; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_94 = 7'h5c == auto_in_a_bits_source ? 6'h2e : _GEN_93; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_95 = 7'h5d == auto_in_a_bits_source ? 6'h2e : _GEN_94; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_96 = 7'h5e == auto_in_a_bits_source ? 6'h2f : _GEN_95; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_97 = 7'h5f == auto_in_a_bits_source ? 6'h2f : _GEN_96; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_98 = 7'h60 == auto_in_a_bits_source ? 6'h30 : _GEN_97; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_99 = 7'h61 == auto_in_a_bits_source ? 6'h30 : _GEN_98; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_100 = 7'h62 == auto_in_a_bits_source ? 6'h31 : _GEN_99; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_101 = 7'h63 == auto_in_a_bits_source ? 6'h31 : _GEN_100; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_102 = 7'h64 == auto_in_a_bits_source ? 6'h32 : _GEN_101; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_103 = 7'h65 == auto_in_a_bits_source ? 6'h32 : _GEN_102; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_104 = 7'h66 == auto_in_a_bits_source ? 6'h33 : _GEN_103; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_105 = 7'h67 == auto_in_a_bits_source ? 6'h33 : _GEN_104; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_106 = 7'h68 == auto_in_a_bits_source ? 6'h34 : _GEN_105; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_107 = 7'h69 == auto_in_a_bits_source ? 6'h34 : _GEN_106; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_108 = 7'h6a == auto_in_a_bits_source ? 6'h35 : _GEN_107; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_109 = 7'h6b == auto_in_a_bits_source ? 6'h35 : _GEN_108; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_110 = 7'h6c == auto_in_a_bits_source ? 6'h36 : _GEN_109; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_111 = 7'h6d == auto_in_a_bits_source ? 6'h36 : _GEN_110; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_112 = 7'h6e == auto_in_a_bits_source ? 6'h37 : _GEN_111; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_113 = 7'h6f == auto_in_a_bits_source ? 6'h37 : _GEN_112; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_114 = 7'h70 == auto_in_a_bits_source ? 6'h38 : _GEN_113; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_115 = 7'h71 == auto_in_a_bits_source ? 6'h38 : _GEN_114; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_116 = 7'h72 == auto_in_a_bits_source ? 6'h39 : _GEN_115; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_117 = 7'h73 == auto_in_a_bits_source ? 6'h39 : _GEN_116; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_118 = 7'h74 == auto_in_a_bits_source ? 6'h3a : _GEN_117; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_119 = 7'h75 == auto_in_a_bits_source ? 6'h3a : _GEN_118; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_120 = 7'h76 == auto_in_a_bits_source ? 6'h3b : _GEN_119; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_121 = 7'h77 == auto_in_a_bits_source ? 6'h3b : _GEN_120; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_122 = 7'h78 == auto_in_a_bits_source ? 6'h3c : _GEN_121; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_123 = 7'h79 == auto_in_a_bits_source ? 6'h3c : _GEN_122; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_124 = 7'h7a == auto_in_a_bits_source ? 6'h3d : _GEN_123; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_125 = 7'h7b == auto_in_a_bits_source ? 6'h3d : _GEN_124; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_126 = 7'h7c == auto_in_a_bits_source ? 6'h3e : _GEN_125; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_127 = 7'h7d == auto_in_a_bits_source ? 6'h3e : _GEN_126; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_128 = 7'h7e == auto_in_a_bits_source ? 6'h3f : _GEN_127; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _GEN_129 = 7'h7f == auto_in_a_bits_source ? 6'h3f : _GEN_128; // @[ToAXI4.scala 165:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292580.4]
  assign _T_962 = 18'h7ff << auto_in_a_bits_size; // @[package.scala 185:77:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292583.4]
  assign _T_963 = _T_962[10:0]; // @[package.scala 185:82:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292584.4]
  assign _T_964 = ~ _T_963; // @[package.scala 185:46:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292585.4]
  assign _T_966 = auto_in_a_bits_size >= 3'h3; // @[ToAXI4.scala 168:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292588.4]
  assign _T_976 = _T_970 & auto_in_a_valid; // @[ToAXI4.scala 178:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292605.4]
  assign _T_977 = _T_957 == 1'h0; // @[ToAXI4.scala 178:61:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292606.4]
  assign _T_978 = _T_977 & _T_933_ready; // @[ToAXI4.scala 178:69:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292607.4]
  assign _T_979 = _T_888 ? _T_978 : 1'h1; // @[ToAXI4.scala 178:51:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292608.4]
  assign _T_980 = _T_976 & _T_979; // @[ToAXI4.scala 178:45:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292609.4]
  assign _T_983 = _T_976 & _T_888; // @[ToAXI4.scala 180:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292613.4]
  assign _T_988 = auto_in_d_ready & auto_out_r_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292621.4]
  assign _T_989 = auto_out_r_bits_last == 1'h0; // @[ToAXI4.scala 188:42:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292623.6]
  assign _T_990 = auto_out_r_valid | _T_987; // @[ToAXI4.scala 190:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292626.4]
  assign _T_991 = _T_990 == 1'h0; // @[ToAXI4.scala 193:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292628.4]
  assign _T_993 = _T_990 ? auto_out_r_valid : auto_out_b_valid; // @[ToAXI4.scala 194:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292631.4]
  assign _T_997 = auto_out_r_bits_resp == 2'h3; // @[ToAXI4.scala 201:39:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292638.4]
  assign _GEN_260 = _T_995 ? _T_997 : _T_999; // @[Reg.scala 12:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292640.4]
  assign _T_1001 = auto_out_r_bits_resp != 2'h0; // @[ToAXI4.scala 202:39:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292644.4]
  assign _T_1002 = auto_out_b_bits_resp != 2'h0; // @[ToAXI4.scala 203:39:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292645.4]
  assign _T_1003 = _T_1001 | _GEN_260; // @[ToAXI4.scala 205:100:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292646.4]
  assign _T_1010 = 64'h1 << _GEN_129; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292671.4]
  assign _T_1012 = _T_1010[0]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292673.4]
  assign _T_1013 = _T_1010[1]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292674.4]
  assign _T_1014 = _T_1010[2]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292675.4]
  assign _T_1015 = _T_1010[3]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292676.4]
  assign _T_1016 = _T_1010[4]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292677.4]
  assign _T_1017 = _T_1010[5]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292678.4]
  assign _T_1018 = _T_1010[6]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292679.4]
  assign _T_1019 = _T_1010[7]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292680.4]
  assign _T_1020 = _T_1010[8]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292681.4]
  assign _T_1021 = _T_1010[9]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292682.4]
  assign _T_1022 = _T_1010[10]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292683.4]
  assign _T_1023 = _T_1010[11]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292684.4]
  assign _T_1024 = _T_1010[12]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292685.4]
  assign _T_1025 = _T_1010[13]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292686.4]
  assign _T_1026 = _T_1010[14]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292687.4]
  assign _T_1027 = _T_1010[15]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292688.4]
  assign _T_1028 = _T_1010[16]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292689.4]
  assign _T_1029 = _T_1010[17]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292690.4]
  assign _T_1030 = _T_1010[18]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292691.4]
  assign _T_1031 = _T_1010[19]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292692.4]
  assign _T_1032 = _T_1010[20]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292693.4]
  assign _T_1033 = _T_1010[21]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292694.4]
  assign _T_1034 = _T_1010[22]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292695.4]
  assign _T_1035 = _T_1010[23]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292696.4]
  assign _T_1036 = _T_1010[24]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292697.4]
  assign _T_1037 = _T_1010[25]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292698.4]
  assign _T_1038 = _T_1010[26]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292699.4]
  assign _T_1039 = _T_1010[27]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292700.4]
  assign _T_1040 = _T_1010[28]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292701.4]
  assign _T_1041 = _T_1010[29]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292702.4]
  assign _T_1042 = _T_1010[30]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292703.4]
  assign _T_1043 = _T_1010[31]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292704.4]
  assign _T_1044 = _T_1010[32]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292705.4]
  assign _T_1045 = _T_1010[33]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292706.4]
  assign _T_1046 = _T_1010[34]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292707.4]
  assign _T_1047 = _T_1010[35]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292708.4]
  assign _T_1048 = _T_1010[36]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292709.4]
  assign _T_1049 = _T_1010[37]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292710.4]
  assign _T_1050 = _T_1010[38]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292711.4]
  assign _T_1051 = _T_1010[39]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292712.4]
  assign _T_1052 = _T_1010[40]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292713.4]
  assign _T_1053 = _T_1010[41]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292714.4]
  assign _T_1054 = _T_1010[42]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292715.4]
  assign _T_1055 = _T_1010[43]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292716.4]
  assign _T_1056 = _T_1010[44]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292717.4]
  assign _T_1057 = _T_1010[45]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292718.4]
  assign _T_1058 = _T_1010[46]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292719.4]
  assign _T_1059 = _T_1010[47]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292720.4]
  assign _T_1060 = _T_1010[48]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292721.4]
  assign _T_1061 = _T_1010[49]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292722.4]
  assign _T_1062 = _T_1010[50]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292723.4]
  assign _T_1063 = _T_1010[51]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292724.4]
  assign _T_1064 = _T_1010[52]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292725.4]
  assign _T_1065 = _T_1010[53]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292726.4]
  assign _T_1066 = _T_1010[54]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292727.4]
  assign _T_1067 = _T_1010[55]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292728.4]
  assign _T_1068 = _T_1010[56]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292729.4]
  assign _T_1069 = _T_1010[57]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292730.4]
  assign _T_1070 = _T_1010[58]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292731.4]
  assign _T_1071 = _T_1010[59]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292732.4]
  assign _T_1072 = _T_1010[60]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292733.4]
  assign _T_1073 = _T_1010[61]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292734.4]
  assign _T_1074 = _T_1010[62]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292735.4]
  assign _T_1075 = _T_1010[63]; // @[ToAXI4.scala 213:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292736.4]
  assign _T_1076 = _T_990 ? auto_out_r_bits_id : auto_out_b_bits_id; // @[ToAXI4.scala 214:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292737.4]
  assign _T_1078 = 64'h1 << _T_1076; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292739.4]
  assign _T_1080 = _T_1078[0]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292741.4]
  assign _T_1081 = _T_1078[1]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292742.4]
  assign _T_1082 = _T_1078[2]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292743.4]
  assign _T_1083 = _T_1078[3]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292744.4]
  assign _T_1084 = _T_1078[4]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292745.4]
  assign _T_1085 = _T_1078[5]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292746.4]
  assign _T_1086 = _T_1078[6]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292747.4]
  assign _T_1087 = _T_1078[7]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292748.4]
  assign _T_1088 = _T_1078[8]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292749.4]
  assign _T_1089 = _T_1078[9]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292750.4]
  assign _T_1090 = _T_1078[10]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292751.4]
  assign _T_1091 = _T_1078[11]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292752.4]
  assign _T_1092 = _T_1078[12]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292753.4]
  assign _T_1093 = _T_1078[13]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292754.4]
  assign _T_1094 = _T_1078[14]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292755.4]
  assign _T_1095 = _T_1078[15]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292756.4]
  assign _T_1096 = _T_1078[16]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292757.4]
  assign _T_1097 = _T_1078[17]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292758.4]
  assign _T_1098 = _T_1078[18]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292759.4]
  assign _T_1099 = _T_1078[19]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292760.4]
  assign _T_1100 = _T_1078[20]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292761.4]
  assign _T_1101 = _T_1078[21]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292762.4]
  assign _T_1102 = _T_1078[22]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292763.4]
  assign _T_1103 = _T_1078[23]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292764.4]
  assign _T_1104 = _T_1078[24]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292765.4]
  assign _T_1105 = _T_1078[25]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292766.4]
  assign _T_1106 = _T_1078[26]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292767.4]
  assign _T_1107 = _T_1078[27]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292768.4]
  assign _T_1108 = _T_1078[28]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292769.4]
  assign _T_1109 = _T_1078[29]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292770.4]
  assign _T_1110 = _T_1078[30]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292771.4]
  assign _T_1111 = _T_1078[31]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292772.4]
  assign _T_1112 = _T_1078[32]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292773.4]
  assign _T_1113 = _T_1078[33]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292774.4]
  assign _T_1114 = _T_1078[34]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292775.4]
  assign _T_1115 = _T_1078[35]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292776.4]
  assign _T_1116 = _T_1078[36]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292777.4]
  assign _T_1117 = _T_1078[37]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292778.4]
  assign _T_1118 = _T_1078[38]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292779.4]
  assign _T_1119 = _T_1078[39]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292780.4]
  assign _T_1120 = _T_1078[40]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292781.4]
  assign _T_1121 = _T_1078[41]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292782.4]
  assign _T_1122 = _T_1078[42]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292783.4]
  assign _T_1123 = _T_1078[43]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292784.4]
  assign _T_1124 = _T_1078[44]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292785.4]
  assign _T_1125 = _T_1078[45]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292786.4]
  assign _T_1126 = _T_1078[46]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292787.4]
  assign _T_1127 = _T_1078[47]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292788.4]
  assign _T_1128 = _T_1078[48]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292789.4]
  assign _T_1129 = _T_1078[49]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292790.4]
  assign _T_1130 = _T_1078[50]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292791.4]
  assign _T_1131 = _T_1078[51]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292792.4]
  assign _T_1132 = _T_1078[52]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292793.4]
  assign _T_1133 = _T_1078[53]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292794.4]
  assign _T_1134 = _T_1078[54]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292795.4]
  assign _T_1135 = _T_1078[55]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292796.4]
  assign _T_1136 = _T_1078[56]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292797.4]
  assign _T_1137 = _T_1078[57]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292798.4]
  assign _T_1138 = _T_1078[58]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292799.4]
  assign _T_1139 = _T_1078[59]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292800.4]
  assign _T_1140 = _T_1078[60]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292801.4]
  assign _T_1141 = _T_1078[61]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292802.4]
  assign _T_1142 = _T_1078[62]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292803.4]
  assign _T_1143 = _T_1078[63]; // @[ToAXI4.scala 214:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292804.4]
  assign _T_1144 = _T_990 ? auto_out_r_bits_last : 1'h1; // @[ToAXI4.scala 215:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292805.4]
  assign _T_1150 = _T_930_ready & _T_980; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292809.4]
  assign _T_1151 = _T_1012 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292810.4]
  assign _T_1152 = _T_1080 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292811.4]
  assign _T_1153 = auto_in_d_ready & _T_993; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292812.4]
  assign _T_1154 = _T_1152 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292813.4]
  assign _T_1156 = _T_1146 + _T_1151; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292815.4]
  assign _T_1157 = _T_1156 - _T_1154; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292816.4]
  assign _T_1158 = $unsigned(_T_1157); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292817.4]
  assign _T_1159 = _T_1158[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292818.4]
  assign _T_1160 = _T_1154 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292820.4]
  assign _T_1162 = _T_1160 | _T_1146; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292822.4]
  assign _T_1164 = _T_1162 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292824.4]
  assign _T_1165 = _T_1164 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292825.4]
  assign _T_1166 = _T_1151 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292830.4]
  assign _T_1167 = _T_1146 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292831.4]
  assign _T_1168 = _T_1166 | _T_1167; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292832.4]
  assign _T_1170 = _T_1168 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292834.4]
  assign _T_1171 = _T_1170 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292835.4]
  assign _T_1182 = _T_1013 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292852.4]
  assign _T_1183 = _T_1081 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292853.4]
  assign _T_1185 = _T_1183 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292855.4]
  assign _T_1187 = _T_1177 + _T_1182; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292857.4]
  assign _T_1188 = _T_1187 - _T_1185; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292858.4]
  assign _T_1189 = $unsigned(_T_1188); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292859.4]
  assign _T_1190 = _T_1189[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292860.4]
  assign _T_1191 = _T_1185 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292862.4]
  assign _T_1193 = _T_1191 | _T_1177; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292864.4]
  assign _T_1195 = _T_1193 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292866.4]
  assign _T_1196 = _T_1195 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292867.4]
  assign _T_1197 = _T_1182 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292872.4]
  assign _T_1198 = _T_1177 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292873.4]
  assign _T_1199 = _T_1197 | _T_1198; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292874.4]
  assign _T_1201 = _T_1199 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292876.4]
  assign _T_1202 = _T_1201 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292877.4]
  assign _T_1213 = _T_1014 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292894.4]
  assign _T_1214 = _T_1082 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292895.4]
  assign _T_1216 = _T_1214 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292897.4]
  assign _T_1218 = _T_1208 + _T_1213; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292899.4]
  assign _T_1219 = _T_1218 - _T_1216; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292900.4]
  assign _T_1220 = $unsigned(_T_1219); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292901.4]
  assign _T_1221 = _T_1220[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292902.4]
  assign _T_1222 = _T_1216 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292904.4]
  assign _T_1224 = _T_1222 | _T_1208; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292906.4]
  assign _T_1226 = _T_1224 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292908.4]
  assign _T_1227 = _T_1226 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292909.4]
  assign _T_1228 = _T_1213 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292914.4]
  assign _T_1229 = _T_1208 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292915.4]
  assign _T_1230 = _T_1228 | _T_1229; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292916.4]
  assign _T_1232 = _T_1230 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292918.4]
  assign _T_1233 = _T_1232 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292919.4]
  assign _T_1244 = _T_1015 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292936.4]
  assign _T_1245 = _T_1083 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292937.4]
  assign _T_1247 = _T_1245 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292939.4]
  assign _T_1249 = _T_1239 + _T_1244; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292941.4]
  assign _T_1250 = _T_1249 - _T_1247; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292942.4]
  assign _T_1251 = $unsigned(_T_1250); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292943.4]
  assign _T_1252 = _T_1251[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292944.4]
  assign _T_1253 = _T_1247 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292946.4]
  assign _T_1255 = _T_1253 | _T_1239; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292948.4]
  assign _T_1257 = _T_1255 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292950.4]
  assign _T_1258 = _T_1257 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292951.4]
  assign _T_1259 = _T_1244 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292956.4]
  assign _T_1260 = _T_1239 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292957.4]
  assign _T_1261 = _T_1259 | _T_1260; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292958.4]
  assign _T_1263 = _T_1261 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292960.4]
  assign _T_1264 = _T_1263 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292961.4]
  assign _T_1275 = _T_1016 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292978.4]
  assign _T_1276 = _T_1084 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292979.4]
  assign _T_1278 = _T_1276 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292981.4]
  assign _T_1280 = _T_1270 + _T_1275; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292983.4]
  assign _T_1281 = _T_1280 - _T_1278; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292984.4]
  assign _T_1282 = $unsigned(_T_1281); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292985.4]
  assign _T_1283 = _T_1282[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292986.4]
  assign _T_1284 = _T_1278 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292988.4]
  assign _T_1286 = _T_1284 | _T_1270; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292990.4]
  assign _T_1288 = _T_1286 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292992.4]
  assign _T_1289 = _T_1288 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292993.4]
  assign _T_1290 = _T_1275 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292998.4]
  assign _T_1291 = _T_1270 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292999.4]
  assign _T_1292 = _T_1290 | _T_1291; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293000.4]
  assign _T_1294 = _T_1292 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293002.4]
  assign _T_1295 = _T_1294 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293003.4]
  assign _T_1306 = _T_1017 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293020.4]
  assign _T_1307 = _T_1085 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293021.4]
  assign _T_1309 = _T_1307 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293023.4]
  assign _T_1311 = _T_1301 + _T_1306; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293025.4]
  assign _T_1312 = _T_1311 - _T_1309; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293026.4]
  assign _T_1313 = $unsigned(_T_1312); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293027.4]
  assign _T_1314 = _T_1313[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293028.4]
  assign _T_1315 = _T_1309 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293030.4]
  assign _T_1317 = _T_1315 | _T_1301; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293032.4]
  assign _T_1319 = _T_1317 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293034.4]
  assign _T_1320 = _T_1319 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293035.4]
  assign _T_1321 = _T_1306 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293040.4]
  assign _T_1322 = _T_1301 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293041.4]
  assign _T_1323 = _T_1321 | _T_1322; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293042.4]
  assign _T_1325 = _T_1323 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293044.4]
  assign _T_1326 = _T_1325 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293045.4]
  assign _T_1337 = _T_1018 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293062.4]
  assign _T_1338 = _T_1086 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293063.4]
  assign _T_1340 = _T_1338 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293065.4]
  assign _T_1342 = _T_1332 + _T_1337; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293067.4]
  assign _T_1343 = _T_1342 - _T_1340; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293068.4]
  assign _T_1344 = $unsigned(_T_1343); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293069.4]
  assign _T_1345 = _T_1344[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293070.4]
  assign _T_1346 = _T_1340 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293072.4]
  assign _T_1348 = _T_1346 | _T_1332; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293074.4]
  assign _T_1350 = _T_1348 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293076.4]
  assign _T_1351 = _T_1350 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293077.4]
  assign _T_1352 = _T_1337 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293082.4]
  assign _T_1353 = _T_1332 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293083.4]
  assign _T_1354 = _T_1352 | _T_1353; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293084.4]
  assign _T_1356 = _T_1354 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293086.4]
  assign _T_1357 = _T_1356 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293087.4]
  assign _T_1368 = _T_1019 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293104.4]
  assign _T_1369 = _T_1087 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293105.4]
  assign _T_1371 = _T_1369 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293107.4]
  assign _T_1373 = _T_1363 + _T_1368; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293109.4]
  assign _T_1374 = _T_1373 - _T_1371; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293110.4]
  assign _T_1375 = $unsigned(_T_1374); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293111.4]
  assign _T_1376 = _T_1375[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293112.4]
  assign _T_1377 = _T_1371 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293114.4]
  assign _T_1379 = _T_1377 | _T_1363; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293116.4]
  assign _T_1381 = _T_1379 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293118.4]
  assign _T_1382 = _T_1381 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293119.4]
  assign _T_1383 = _T_1368 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293124.4]
  assign _T_1384 = _T_1363 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293125.4]
  assign _T_1385 = _T_1383 | _T_1384; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293126.4]
  assign _T_1387 = _T_1385 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293128.4]
  assign _T_1388 = _T_1387 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293129.4]
  assign _T_1399 = _T_1020 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293146.4]
  assign _T_1400 = _T_1088 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293147.4]
  assign _T_1402 = _T_1400 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293149.4]
  assign _T_1404 = _T_1394 + _T_1399; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293151.4]
  assign _T_1405 = _T_1404 - _T_1402; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293152.4]
  assign _T_1406 = $unsigned(_T_1405); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293153.4]
  assign _T_1407 = _T_1406[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293154.4]
  assign _T_1408 = _T_1402 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293156.4]
  assign _T_1410 = _T_1408 | _T_1394; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293158.4]
  assign _T_1412 = _T_1410 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293160.4]
  assign _T_1413 = _T_1412 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293161.4]
  assign _T_1414 = _T_1399 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293166.4]
  assign _T_1415 = _T_1394 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293167.4]
  assign _T_1416 = _T_1414 | _T_1415; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293168.4]
  assign _T_1418 = _T_1416 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293170.4]
  assign _T_1419 = _T_1418 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293171.4]
  assign _T_1430 = _T_1021 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293188.4]
  assign _T_1431 = _T_1089 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293189.4]
  assign _T_1433 = _T_1431 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293191.4]
  assign _T_1435 = _T_1425 + _T_1430; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293193.4]
  assign _T_1436 = _T_1435 - _T_1433; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293194.4]
  assign _T_1437 = $unsigned(_T_1436); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293195.4]
  assign _T_1438 = _T_1437[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293196.4]
  assign _T_1439 = _T_1433 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293198.4]
  assign _T_1441 = _T_1439 | _T_1425; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293200.4]
  assign _T_1443 = _T_1441 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293202.4]
  assign _T_1444 = _T_1443 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293203.4]
  assign _T_1445 = _T_1430 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293208.4]
  assign _T_1446 = _T_1425 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293209.4]
  assign _T_1447 = _T_1445 | _T_1446; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293210.4]
  assign _T_1449 = _T_1447 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293212.4]
  assign _T_1450 = _T_1449 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293213.4]
  assign _T_1461 = _T_1022 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293230.4]
  assign _T_1462 = _T_1090 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293231.4]
  assign _T_1464 = _T_1462 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293233.4]
  assign _T_1466 = _T_1456 + _T_1461; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293235.4]
  assign _T_1467 = _T_1466 - _T_1464; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293236.4]
  assign _T_1468 = $unsigned(_T_1467); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293237.4]
  assign _T_1469 = _T_1468[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293238.4]
  assign _T_1470 = _T_1464 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293240.4]
  assign _T_1472 = _T_1470 | _T_1456; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293242.4]
  assign _T_1474 = _T_1472 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293244.4]
  assign _T_1475 = _T_1474 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293245.4]
  assign _T_1476 = _T_1461 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293250.4]
  assign _T_1477 = _T_1456 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293251.4]
  assign _T_1478 = _T_1476 | _T_1477; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293252.4]
  assign _T_1480 = _T_1478 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293254.4]
  assign _T_1481 = _T_1480 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293255.4]
  assign _T_1492 = _T_1023 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293272.4]
  assign _T_1493 = _T_1091 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293273.4]
  assign _T_1495 = _T_1493 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293275.4]
  assign _T_1497 = _T_1487 + _T_1492; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293277.4]
  assign _T_1498 = _T_1497 - _T_1495; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293278.4]
  assign _T_1499 = $unsigned(_T_1498); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293279.4]
  assign _T_1500 = _T_1499[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293280.4]
  assign _T_1501 = _T_1495 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293282.4]
  assign _T_1503 = _T_1501 | _T_1487; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293284.4]
  assign _T_1505 = _T_1503 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293286.4]
  assign _T_1506 = _T_1505 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293287.4]
  assign _T_1507 = _T_1492 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293292.4]
  assign _T_1508 = _T_1487 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293293.4]
  assign _T_1509 = _T_1507 | _T_1508; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293294.4]
  assign _T_1511 = _T_1509 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293296.4]
  assign _T_1512 = _T_1511 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293297.4]
  assign _T_1523 = _T_1024 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293314.4]
  assign _T_1524 = _T_1092 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293315.4]
  assign _T_1526 = _T_1524 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293317.4]
  assign _T_1528 = _T_1518 + _T_1523; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293319.4]
  assign _T_1529 = _T_1528 - _T_1526; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293320.4]
  assign _T_1530 = $unsigned(_T_1529); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293321.4]
  assign _T_1531 = _T_1530[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293322.4]
  assign _T_1532 = _T_1526 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293324.4]
  assign _T_1534 = _T_1532 | _T_1518; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293326.4]
  assign _T_1536 = _T_1534 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293328.4]
  assign _T_1537 = _T_1536 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293329.4]
  assign _T_1538 = _T_1523 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293334.4]
  assign _T_1539 = _T_1518 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293335.4]
  assign _T_1540 = _T_1538 | _T_1539; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293336.4]
  assign _T_1542 = _T_1540 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293338.4]
  assign _T_1543 = _T_1542 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293339.4]
  assign _T_1554 = _T_1025 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293356.4]
  assign _T_1555 = _T_1093 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293357.4]
  assign _T_1557 = _T_1555 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293359.4]
  assign _T_1559 = _T_1549 + _T_1554; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293361.4]
  assign _T_1560 = _T_1559 - _T_1557; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293362.4]
  assign _T_1561 = $unsigned(_T_1560); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293363.4]
  assign _T_1562 = _T_1561[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293364.4]
  assign _T_1563 = _T_1557 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293366.4]
  assign _T_1565 = _T_1563 | _T_1549; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293368.4]
  assign _T_1567 = _T_1565 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293370.4]
  assign _T_1568 = _T_1567 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293371.4]
  assign _T_1569 = _T_1554 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293376.4]
  assign _T_1570 = _T_1549 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293377.4]
  assign _T_1571 = _T_1569 | _T_1570; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293378.4]
  assign _T_1573 = _T_1571 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293380.4]
  assign _T_1574 = _T_1573 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293381.4]
  assign _T_1585 = _T_1026 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293398.4]
  assign _T_1586 = _T_1094 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293399.4]
  assign _T_1588 = _T_1586 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293401.4]
  assign _T_1590 = _T_1580 + _T_1585; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293403.4]
  assign _T_1591 = _T_1590 - _T_1588; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293404.4]
  assign _T_1592 = $unsigned(_T_1591); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293405.4]
  assign _T_1593 = _T_1592[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293406.4]
  assign _T_1594 = _T_1588 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293408.4]
  assign _T_1596 = _T_1594 | _T_1580; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293410.4]
  assign _T_1598 = _T_1596 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293412.4]
  assign _T_1599 = _T_1598 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293413.4]
  assign _T_1600 = _T_1585 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293418.4]
  assign _T_1601 = _T_1580 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293419.4]
  assign _T_1602 = _T_1600 | _T_1601; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293420.4]
  assign _T_1604 = _T_1602 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293422.4]
  assign _T_1605 = _T_1604 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293423.4]
  assign _T_1616 = _T_1027 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293440.4]
  assign _T_1617 = _T_1095 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293441.4]
  assign _T_1619 = _T_1617 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293443.4]
  assign _T_1621 = _T_1611 + _T_1616; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293445.4]
  assign _T_1622 = _T_1621 - _T_1619; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293446.4]
  assign _T_1623 = $unsigned(_T_1622); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293447.4]
  assign _T_1624 = _T_1623[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293448.4]
  assign _T_1625 = _T_1619 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293450.4]
  assign _T_1627 = _T_1625 | _T_1611; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293452.4]
  assign _T_1629 = _T_1627 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293454.4]
  assign _T_1630 = _T_1629 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293455.4]
  assign _T_1631 = _T_1616 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293460.4]
  assign _T_1632 = _T_1611 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293461.4]
  assign _T_1633 = _T_1631 | _T_1632; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293462.4]
  assign _T_1635 = _T_1633 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293464.4]
  assign _T_1636 = _T_1635 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293465.4]
  assign _T_1647 = _T_1028 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293482.4]
  assign _T_1648 = _T_1096 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293483.4]
  assign _T_1650 = _T_1648 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293485.4]
  assign _T_1652 = _T_1642 + _T_1647; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293487.4]
  assign _T_1653 = _T_1652 - _T_1650; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293488.4]
  assign _T_1654 = $unsigned(_T_1653); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293489.4]
  assign _T_1655 = _T_1654[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293490.4]
  assign _T_1656 = _T_1650 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293492.4]
  assign _T_1658 = _T_1656 | _T_1642; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293494.4]
  assign _T_1660 = _T_1658 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293496.4]
  assign _T_1661 = _T_1660 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293497.4]
  assign _T_1662 = _T_1647 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293502.4]
  assign _T_1663 = _T_1642 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293503.4]
  assign _T_1664 = _T_1662 | _T_1663; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293504.4]
  assign _T_1666 = _T_1664 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293506.4]
  assign _T_1667 = _T_1666 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293507.4]
  assign _T_1678 = _T_1029 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293524.4]
  assign _T_1679 = _T_1097 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293525.4]
  assign _T_1681 = _T_1679 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293527.4]
  assign _T_1683 = _T_1673 + _T_1678; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293529.4]
  assign _T_1684 = _T_1683 - _T_1681; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293530.4]
  assign _T_1685 = $unsigned(_T_1684); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293531.4]
  assign _T_1686 = _T_1685[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293532.4]
  assign _T_1687 = _T_1681 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293534.4]
  assign _T_1689 = _T_1687 | _T_1673; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293536.4]
  assign _T_1691 = _T_1689 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293538.4]
  assign _T_1692 = _T_1691 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293539.4]
  assign _T_1693 = _T_1678 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293544.4]
  assign _T_1694 = _T_1673 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293545.4]
  assign _T_1695 = _T_1693 | _T_1694; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293546.4]
  assign _T_1697 = _T_1695 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293548.4]
  assign _T_1698 = _T_1697 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293549.4]
  assign _T_1709 = _T_1030 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293566.4]
  assign _T_1710 = _T_1098 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293567.4]
  assign _T_1712 = _T_1710 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293569.4]
  assign _T_1714 = _T_1704 + _T_1709; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293571.4]
  assign _T_1715 = _T_1714 - _T_1712; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293572.4]
  assign _T_1716 = $unsigned(_T_1715); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293573.4]
  assign _T_1717 = _T_1716[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293574.4]
  assign _T_1718 = _T_1712 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293576.4]
  assign _T_1720 = _T_1718 | _T_1704; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293578.4]
  assign _T_1722 = _T_1720 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293580.4]
  assign _T_1723 = _T_1722 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293581.4]
  assign _T_1724 = _T_1709 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293586.4]
  assign _T_1725 = _T_1704 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293587.4]
  assign _T_1726 = _T_1724 | _T_1725; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293588.4]
  assign _T_1728 = _T_1726 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293590.4]
  assign _T_1729 = _T_1728 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293591.4]
  assign _T_1740 = _T_1031 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293608.4]
  assign _T_1741 = _T_1099 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293609.4]
  assign _T_1743 = _T_1741 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293611.4]
  assign _T_1745 = _T_1735 + _T_1740; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293613.4]
  assign _T_1746 = _T_1745 - _T_1743; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293614.4]
  assign _T_1747 = $unsigned(_T_1746); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293615.4]
  assign _T_1748 = _T_1747[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293616.4]
  assign _T_1749 = _T_1743 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293618.4]
  assign _T_1751 = _T_1749 | _T_1735; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293620.4]
  assign _T_1753 = _T_1751 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293622.4]
  assign _T_1754 = _T_1753 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293623.4]
  assign _T_1755 = _T_1740 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293628.4]
  assign _T_1756 = _T_1735 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293629.4]
  assign _T_1757 = _T_1755 | _T_1756; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293630.4]
  assign _T_1759 = _T_1757 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293632.4]
  assign _T_1760 = _T_1759 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293633.4]
  assign _T_1771 = _T_1032 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293650.4]
  assign _T_1772 = _T_1100 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293651.4]
  assign _T_1774 = _T_1772 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293653.4]
  assign _T_1776 = _T_1766 + _T_1771; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293655.4]
  assign _T_1777 = _T_1776 - _T_1774; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293656.4]
  assign _T_1778 = $unsigned(_T_1777); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293657.4]
  assign _T_1779 = _T_1778[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293658.4]
  assign _T_1780 = _T_1774 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293660.4]
  assign _T_1782 = _T_1780 | _T_1766; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293662.4]
  assign _T_1784 = _T_1782 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293664.4]
  assign _T_1785 = _T_1784 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293665.4]
  assign _T_1786 = _T_1771 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293670.4]
  assign _T_1787 = _T_1766 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293671.4]
  assign _T_1788 = _T_1786 | _T_1787; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293672.4]
  assign _T_1790 = _T_1788 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293674.4]
  assign _T_1791 = _T_1790 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293675.4]
  assign _T_1802 = _T_1033 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293692.4]
  assign _T_1803 = _T_1101 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293693.4]
  assign _T_1805 = _T_1803 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293695.4]
  assign _T_1807 = _T_1797 + _T_1802; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293697.4]
  assign _T_1808 = _T_1807 - _T_1805; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293698.4]
  assign _T_1809 = $unsigned(_T_1808); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293699.4]
  assign _T_1810 = _T_1809[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293700.4]
  assign _T_1811 = _T_1805 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293702.4]
  assign _T_1813 = _T_1811 | _T_1797; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293704.4]
  assign _T_1815 = _T_1813 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293706.4]
  assign _T_1816 = _T_1815 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293707.4]
  assign _T_1817 = _T_1802 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293712.4]
  assign _T_1818 = _T_1797 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293713.4]
  assign _T_1819 = _T_1817 | _T_1818; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293714.4]
  assign _T_1821 = _T_1819 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293716.4]
  assign _T_1822 = _T_1821 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293717.4]
  assign _T_1833 = _T_1034 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293734.4]
  assign _T_1834 = _T_1102 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293735.4]
  assign _T_1836 = _T_1834 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293737.4]
  assign _T_1838 = _T_1828 + _T_1833; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293739.4]
  assign _T_1839 = _T_1838 - _T_1836; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293740.4]
  assign _T_1840 = $unsigned(_T_1839); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293741.4]
  assign _T_1841 = _T_1840[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293742.4]
  assign _T_1842 = _T_1836 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293744.4]
  assign _T_1844 = _T_1842 | _T_1828; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293746.4]
  assign _T_1846 = _T_1844 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293748.4]
  assign _T_1847 = _T_1846 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293749.4]
  assign _T_1848 = _T_1833 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293754.4]
  assign _T_1849 = _T_1828 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293755.4]
  assign _T_1850 = _T_1848 | _T_1849; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293756.4]
  assign _T_1852 = _T_1850 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293758.4]
  assign _T_1853 = _T_1852 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293759.4]
  assign _T_1864 = _T_1035 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293776.4]
  assign _T_1865 = _T_1103 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293777.4]
  assign _T_1867 = _T_1865 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293779.4]
  assign _T_1869 = _T_1859 + _T_1864; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293781.4]
  assign _T_1870 = _T_1869 - _T_1867; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293782.4]
  assign _T_1871 = $unsigned(_T_1870); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293783.4]
  assign _T_1872 = _T_1871[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293784.4]
  assign _T_1873 = _T_1867 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293786.4]
  assign _T_1875 = _T_1873 | _T_1859; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293788.4]
  assign _T_1877 = _T_1875 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293790.4]
  assign _T_1878 = _T_1877 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293791.4]
  assign _T_1879 = _T_1864 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293796.4]
  assign _T_1880 = _T_1859 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293797.4]
  assign _T_1881 = _T_1879 | _T_1880; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293798.4]
  assign _T_1883 = _T_1881 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293800.4]
  assign _T_1884 = _T_1883 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293801.4]
  assign _T_1895 = _T_1036 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293818.4]
  assign _T_1896 = _T_1104 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293819.4]
  assign _T_1898 = _T_1896 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293821.4]
  assign _T_1900 = _T_1890 + _T_1895; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293823.4]
  assign _T_1901 = _T_1900 - _T_1898; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293824.4]
  assign _T_1902 = $unsigned(_T_1901); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293825.4]
  assign _T_1903 = _T_1902[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293826.4]
  assign _T_1904 = _T_1898 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293828.4]
  assign _T_1906 = _T_1904 | _T_1890; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293830.4]
  assign _T_1908 = _T_1906 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293832.4]
  assign _T_1909 = _T_1908 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293833.4]
  assign _T_1910 = _T_1895 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293838.4]
  assign _T_1911 = _T_1890 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293839.4]
  assign _T_1912 = _T_1910 | _T_1911; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293840.4]
  assign _T_1914 = _T_1912 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293842.4]
  assign _T_1915 = _T_1914 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293843.4]
  assign _T_1926 = _T_1037 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293860.4]
  assign _T_1927 = _T_1105 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293861.4]
  assign _T_1929 = _T_1927 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293863.4]
  assign _T_1931 = _T_1921 + _T_1926; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293865.4]
  assign _T_1932 = _T_1931 - _T_1929; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293866.4]
  assign _T_1933 = $unsigned(_T_1932); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293867.4]
  assign _T_1934 = _T_1933[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293868.4]
  assign _T_1935 = _T_1929 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293870.4]
  assign _T_1937 = _T_1935 | _T_1921; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293872.4]
  assign _T_1939 = _T_1937 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293874.4]
  assign _T_1940 = _T_1939 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293875.4]
  assign _T_1941 = _T_1926 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293880.4]
  assign _T_1942 = _T_1921 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293881.4]
  assign _T_1943 = _T_1941 | _T_1942; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293882.4]
  assign _T_1945 = _T_1943 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293884.4]
  assign _T_1946 = _T_1945 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293885.4]
  assign _T_1957 = _T_1038 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293902.4]
  assign _T_1958 = _T_1106 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293903.4]
  assign _T_1960 = _T_1958 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293905.4]
  assign _T_1962 = _T_1952 + _T_1957; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293907.4]
  assign _T_1963 = _T_1962 - _T_1960; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293908.4]
  assign _T_1964 = $unsigned(_T_1963); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293909.4]
  assign _T_1965 = _T_1964[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293910.4]
  assign _T_1966 = _T_1960 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293912.4]
  assign _T_1968 = _T_1966 | _T_1952; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293914.4]
  assign _T_1970 = _T_1968 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293916.4]
  assign _T_1971 = _T_1970 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293917.4]
  assign _T_1972 = _T_1957 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293922.4]
  assign _T_1973 = _T_1952 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293923.4]
  assign _T_1974 = _T_1972 | _T_1973; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293924.4]
  assign _T_1976 = _T_1974 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293926.4]
  assign _T_1977 = _T_1976 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293927.4]
  assign _T_1988 = _T_1039 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293944.4]
  assign _T_1989 = _T_1107 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293945.4]
  assign _T_1991 = _T_1989 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293947.4]
  assign _T_1993 = _T_1983 + _T_1988; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293949.4]
  assign _T_1994 = _T_1993 - _T_1991; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293950.4]
  assign _T_1995 = $unsigned(_T_1994); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293951.4]
  assign _T_1996 = _T_1995[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293952.4]
  assign _T_1997 = _T_1991 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293954.4]
  assign _T_1999 = _T_1997 | _T_1983; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293956.4]
  assign _T_2001 = _T_1999 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293958.4]
  assign _T_2002 = _T_2001 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293959.4]
  assign _T_2003 = _T_1988 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293964.4]
  assign _T_2004 = _T_1983 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293965.4]
  assign _T_2005 = _T_2003 | _T_2004; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293966.4]
  assign _T_2007 = _T_2005 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293968.4]
  assign _T_2008 = _T_2007 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293969.4]
  assign _T_2019 = _T_1040 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293986.4]
  assign _T_2020 = _T_1108 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293987.4]
  assign _T_2022 = _T_2020 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293989.4]
  assign _T_2024 = _T_2014 + _T_2019; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293991.4]
  assign _T_2025 = _T_2024 - _T_2022; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293992.4]
  assign _T_2026 = $unsigned(_T_2025); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293993.4]
  assign _T_2027 = _T_2026[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293994.4]
  assign _T_2028 = _T_2022 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293996.4]
  assign _T_2030 = _T_2028 | _T_2014; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293998.4]
  assign _T_2032 = _T_2030 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294000.4]
  assign _T_2033 = _T_2032 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294001.4]
  assign _T_2034 = _T_2019 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294006.4]
  assign _T_2035 = _T_2014 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294007.4]
  assign _T_2036 = _T_2034 | _T_2035; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294008.4]
  assign _T_2038 = _T_2036 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294010.4]
  assign _T_2039 = _T_2038 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294011.4]
  assign _T_2050 = _T_1041 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294028.4]
  assign _T_2051 = _T_1109 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294029.4]
  assign _T_2053 = _T_2051 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294031.4]
  assign _T_2055 = _T_2045 + _T_2050; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294033.4]
  assign _T_2056 = _T_2055 - _T_2053; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294034.4]
  assign _T_2057 = $unsigned(_T_2056); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294035.4]
  assign _T_2058 = _T_2057[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294036.4]
  assign _T_2059 = _T_2053 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294038.4]
  assign _T_2061 = _T_2059 | _T_2045; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294040.4]
  assign _T_2063 = _T_2061 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294042.4]
  assign _T_2064 = _T_2063 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294043.4]
  assign _T_2065 = _T_2050 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294048.4]
  assign _T_2066 = _T_2045 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294049.4]
  assign _T_2067 = _T_2065 | _T_2066; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294050.4]
  assign _T_2069 = _T_2067 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294052.4]
  assign _T_2070 = _T_2069 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294053.4]
  assign _T_2081 = _T_1042 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294070.4]
  assign _T_2082 = _T_1110 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294071.4]
  assign _T_2084 = _T_2082 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294073.4]
  assign _T_2086 = _T_2076 + _T_2081; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294075.4]
  assign _T_2087 = _T_2086 - _T_2084; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294076.4]
  assign _T_2088 = $unsigned(_T_2087); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294077.4]
  assign _T_2089 = _T_2088[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294078.4]
  assign _T_2090 = _T_2084 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294080.4]
  assign _T_2092 = _T_2090 | _T_2076; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294082.4]
  assign _T_2094 = _T_2092 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294084.4]
  assign _T_2095 = _T_2094 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294085.4]
  assign _T_2096 = _T_2081 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294090.4]
  assign _T_2097 = _T_2076 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294091.4]
  assign _T_2098 = _T_2096 | _T_2097; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294092.4]
  assign _T_2100 = _T_2098 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294094.4]
  assign _T_2101 = _T_2100 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294095.4]
  assign _T_2112 = _T_1043 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294112.4]
  assign _T_2113 = _T_1111 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294113.4]
  assign _T_2115 = _T_2113 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294115.4]
  assign _T_2117 = _T_2107 + _T_2112; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294117.4]
  assign _T_2118 = _T_2117 - _T_2115; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294118.4]
  assign _T_2119 = $unsigned(_T_2118); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294119.4]
  assign _T_2120 = _T_2119[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294120.4]
  assign _T_2121 = _T_2115 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294122.4]
  assign _T_2123 = _T_2121 | _T_2107; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294124.4]
  assign _T_2125 = _T_2123 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294126.4]
  assign _T_2126 = _T_2125 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294127.4]
  assign _T_2127 = _T_2112 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294132.4]
  assign _T_2128 = _T_2107 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294133.4]
  assign _T_2129 = _T_2127 | _T_2128; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294134.4]
  assign _T_2131 = _T_2129 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294136.4]
  assign _T_2132 = _T_2131 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294137.4]
  assign _T_2143 = _T_1044 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294154.4]
  assign _T_2144 = _T_1112 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294155.4]
  assign _T_2146 = _T_2144 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294157.4]
  assign _T_2148 = _T_2138 + _T_2143; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294159.4]
  assign _T_2149 = _T_2148 - _T_2146; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294160.4]
  assign _T_2150 = $unsigned(_T_2149); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294161.4]
  assign _T_2151 = _T_2150[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294162.4]
  assign _T_2152 = _T_2146 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294164.4]
  assign _T_2154 = _T_2152 | _T_2138; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294166.4]
  assign _T_2156 = _T_2154 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294168.4]
  assign _T_2157 = _T_2156 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294169.4]
  assign _T_2158 = _T_2143 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294174.4]
  assign _T_2159 = _T_2138 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294175.4]
  assign _T_2160 = _T_2158 | _T_2159; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294176.4]
  assign _T_2162 = _T_2160 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294178.4]
  assign _T_2163 = _T_2162 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294179.4]
  assign _T_2174 = _T_1045 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294196.4]
  assign _T_2175 = _T_1113 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294197.4]
  assign _T_2177 = _T_2175 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294199.4]
  assign _T_2179 = _T_2169 + _T_2174; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294201.4]
  assign _T_2180 = _T_2179 - _T_2177; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294202.4]
  assign _T_2181 = $unsigned(_T_2180); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294203.4]
  assign _T_2182 = _T_2181[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294204.4]
  assign _T_2183 = _T_2177 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294206.4]
  assign _T_2185 = _T_2183 | _T_2169; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294208.4]
  assign _T_2187 = _T_2185 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294210.4]
  assign _T_2188 = _T_2187 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294211.4]
  assign _T_2189 = _T_2174 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294216.4]
  assign _T_2190 = _T_2169 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294217.4]
  assign _T_2191 = _T_2189 | _T_2190; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294218.4]
  assign _T_2193 = _T_2191 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294220.4]
  assign _T_2194 = _T_2193 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294221.4]
  assign _T_2205 = _T_1046 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294238.4]
  assign _T_2206 = _T_1114 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294239.4]
  assign _T_2208 = _T_2206 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294241.4]
  assign _T_2210 = _T_2200 + _T_2205; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294243.4]
  assign _T_2211 = _T_2210 - _T_2208; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294244.4]
  assign _T_2212 = $unsigned(_T_2211); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294245.4]
  assign _T_2213 = _T_2212[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294246.4]
  assign _T_2214 = _T_2208 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294248.4]
  assign _T_2216 = _T_2214 | _T_2200; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294250.4]
  assign _T_2218 = _T_2216 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294252.4]
  assign _T_2219 = _T_2218 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294253.4]
  assign _T_2220 = _T_2205 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294258.4]
  assign _T_2221 = _T_2200 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294259.4]
  assign _T_2222 = _T_2220 | _T_2221; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294260.4]
  assign _T_2224 = _T_2222 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294262.4]
  assign _T_2225 = _T_2224 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294263.4]
  assign _T_2236 = _T_1047 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294280.4]
  assign _T_2237 = _T_1115 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294281.4]
  assign _T_2239 = _T_2237 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294283.4]
  assign _T_2241 = _T_2231 + _T_2236; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294285.4]
  assign _T_2242 = _T_2241 - _T_2239; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294286.4]
  assign _T_2243 = $unsigned(_T_2242); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294287.4]
  assign _T_2244 = _T_2243[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294288.4]
  assign _T_2245 = _T_2239 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294290.4]
  assign _T_2247 = _T_2245 | _T_2231; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294292.4]
  assign _T_2249 = _T_2247 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294294.4]
  assign _T_2250 = _T_2249 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294295.4]
  assign _T_2251 = _T_2236 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294300.4]
  assign _T_2252 = _T_2231 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294301.4]
  assign _T_2253 = _T_2251 | _T_2252; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294302.4]
  assign _T_2255 = _T_2253 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294304.4]
  assign _T_2256 = _T_2255 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294305.4]
  assign _T_2267 = _T_1048 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294322.4]
  assign _T_2268 = _T_1116 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294323.4]
  assign _T_2270 = _T_2268 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294325.4]
  assign _T_2272 = _T_2262 + _T_2267; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294327.4]
  assign _T_2273 = _T_2272 - _T_2270; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294328.4]
  assign _T_2274 = $unsigned(_T_2273); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294329.4]
  assign _T_2275 = _T_2274[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294330.4]
  assign _T_2276 = _T_2270 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294332.4]
  assign _T_2278 = _T_2276 | _T_2262; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294334.4]
  assign _T_2280 = _T_2278 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294336.4]
  assign _T_2281 = _T_2280 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294337.4]
  assign _T_2282 = _T_2267 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294342.4]
  assign _T_2283 = _T_2262 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294343.4]
  assign _T_2284 = _T_2282 | _T_2283; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294344.4]
  assign _T_2286 = _T_2284 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294346.4]
  assign _T_2287 = _T_2286 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294347.4]
  assign _T_2298 = _T_1049 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294364.4]
  assign _T_2299 = _T_1117 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294365.4]
  assign _T_2301 = _T_2299 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294367.4]
  assign _T_2303 = _T_2293 + _T_2298; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294369.4]
  assign _T_2304 = _T_2303 - _T_2301; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294370.4]
  assign _T_2305 = $unsigned(_T_2304); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294371.4]
  assign _T_2306 = _T_2305[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294372.4]
  assign _T_2307 = _T_2301 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294374.4]
  assign _T_2309 = _T_2307 | _T_2293; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294376.4]
  assign _T_2311 = _T_2309 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294378.4]
  assign _T_2312 = _T_2311 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294379.4]
  assign _T_2313 = _T_2298 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294384.4]
  assign _T_2314 = _T_2293 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294385.4]
  assign _T_2315 = _T_2313 | _T_2314; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294386.4]
  assign _T_2317 = _T_2315 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294388.4]
  assign _T_2318 = _T_2317 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294389.4]
  assign _T_2329 = _T_1050 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294406.4]
  assign _T_2330 = _T_1118 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294407.4]
  assign _T_2332 = _T_2330 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294409.4]
  assign _T_2334 = _T_2324 + _T_2329; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294411.4]
  assign _T_2335 = _T_2334 - _T_2332; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294412.4]
  assign _T_2336 = $unsigned(_T_2335); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294413.4]
  assign _T_2337 = _T_2336[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294414.4]
  assign _T_2338 = _T_2332 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294416.4]
  assign _T_2340 = _T_2338 | _T_2324; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294418.4]
  assign _T_2342 = _T_2340 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294420.4]
  assign _T_2343 = _T_2342 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294421.4]
  assign _T_2344 = _T_2329 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294426.4]
  assign _T_2345 = _T_2324 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294427.4]
  assign _T_2346 = _T_2344 | _T_2345; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294428.4]
  assign _T_2348 = _T_2346 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294430.4]
  assign _T_2349 = _T_2348 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294431.4]
  assign _T_2360 = _T_1051 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294448.4]
  assign _T_2361 = _T_1119 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294449.4]
  assign _T_2363 = _T_2361 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294451.4]
  assign _T_2365 = _T_2355 + _T_2360; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294453.4]
  assign _T_2366 = _T_2365 - _T_2363; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294454.4]
  assign _T_2367 = $unsigned(_T_2366); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294455.4]
  assign _T_2368 = _T_2367[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294456.4]
  assign _T_2369 = _T_2363 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294458.4]
  assign _T_2371 = _T_2369 | _T_2355; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294460.4]
  assign _T_2373 = _T_2371 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294462.4]
  assign _T_2374 = _T_2373 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294463.4]
  assign _T_2375 = _T_2360 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294468.4]
  assign _T_2376 = _T_2355 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294469.4]
  assign _T_2377 = _T_2375 | _T_2376; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294470.4]
  assign _T_2379 = _T_2377 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294472.4]
  assign _T_2380 = _T_2379 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294473.4]
  assign _T_2391 = _T_1052 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294490.4]
  assign _T_2392 = _T_1120 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294491.4]
  assign _T_2394 = _T_2392 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294493.4]
  assign _T_2396 = _T_2386 + _T_2391; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294495.4]
  assign _T_2397 = _T_2396 - _T_2394; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294496.4]
  assign _T_2398 = $unsigned(_T_2397); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294497.4]
  assign _T_2399 = _T_2398[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294498.4]
  assign _T_2400 = _T_2394 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294500.4]
  assign _T_2402 = _T_2400 | _T_2386; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294502.4]
  assign _T_2404 = _T_2402 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294504.4]
  assign _T_2405 = _T_2404 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294505.4]
  assign _T_2406 = _T_2391 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294510.4]
  assign _T_2407 = _T_2386 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294511.4]
  assign _T_2408 = _T_2406 | _T_2407; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294512.4]
  assign _T_2410 = _T_2408 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294514.4]
  assign _T_2411 = _T_2410 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294515.4]
  assign _T_2422 = _T_1053 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294532.4]
  assign _T_2423 = _T_1121 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294533.4]
  assign _T_2425 = _T_2423 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294535.4]
  assign _T_2427 = _T_2417 + _T_2422; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294537.4]
  assign _T_2428 = _T_2427 - _T_2425; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294538.4]
  assign _T_2429 = $unsigned(_T_2428); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294539.4]
  assign _T_2430 = _T_2429[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294540.4]
  assign _T_2431 = _T_2425 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294542.4]
  assign _T_2433 = _T_2431 | _T_2417; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294544.4]
  assign _T_2435 = _T_2433 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294546.4]
  assign _T_2436 = _T_2435 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294547.4]
  assign _T_2437 = _T_2422 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294552.4]
  assign _T_2438 = _T_2417 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294553.4]
  assign _T_2439 = _T_2437 | _T_2438; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294554.4]
  assign _T_2441 = _T_2439 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294556.4]
  assign _T_2442 = _T_2441 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294557.4]
  assign _T_2453 = _T_1054 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294574.4]
  assign _T_2454 = _T_1122 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294575.4]
  assign _T_2456 = _T_2454 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294577.4]
  assign _T_2458 = _T_2448 + _T_2453; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294579.4]
  assign _T_2459 = _T_2458 - _T_2456; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294580.4]
  assign _T_2460 = $unsigned(_T_2459); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294581.4]
  assign _T_2461 = _T_2460[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294582.4]
  assign _T_2462 = _T_2456 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294584.4]
  assign _T_2464 = _T_2462 | _T_2448; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294586.4]
  assign _T_2466 = _T_2464 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294588.4]
  assign _T_2467 = _T_2466 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294589.4]
  assign _T_2468 = _T_2453 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294594.4]
  assign _T_2469 = _T_2448 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294595.4]
  assign _T_2470 = _T_2468 | _T_2469; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294596.4]
  assign _T_2472 = _T_2470 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294598.4]
  assign _T_2473 = _T_2472 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294599.4]
  assign _T_2484 = _T_1055 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294616.4]
  assign _T_2485 = _T_1123 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294617.4]
  assign _T_2487 = _T_2485 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294619.4]
  assign _T_2489 = _T_2479 + _T_2484; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294621.4]
  assign _T_2490 = _T_2489 - _T_2487; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294622.4]
  assign _T_2491 = $unsigned(_T_2490); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294623.4]
  assign _T_2492 = _T_2491[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294624.4]
  assign _T_2493 = _T_2487 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294626.4]
  assign _T_2495 = _T_2493 | _T_2479; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294628.4]
  assign _T_2497 = _T_2495 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294630.4]
  assign _T_2498 = _T_2497 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294631.4]
  assign _T_2499 = _T_2484 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294636.4]
  assign _T_2500 = _T_2479 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294637.4]
  assign _T_2501 = _T_2499 | _T_2500; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294638.4]
  assign _T_2503 = _T_2501 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294640.4]
  assign _T_2504 = _T_2503 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294641.4]
  assign _T_2515 = _T_1056 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294658.4]
  assign _T_2516 = _T_1124 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294659.4]
  assign _T_2518 = _T_2516 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294661.4]
  assign _T_2520 = _T_2510 + _T_2515; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294663.4]
  assign _T_2521 = _T_2520 - _T_2518; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294664.4]
  assign _T_2522 = $unsigned(_T_2521); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294665.4]
  assign _T_2523 = _T_2522[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294666.4]
  assign _T_2524 = _T_2518 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294668.4]
  assign _T_2526 = _T_2524 | _T_2510; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294670.4]
  assign _T_2528 = _T_2526 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294672.4]
  assign _T_2529 = _T_2528 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294673.4]
  assign _T_2530 = _T_2515 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294678.4]
  assign _T_2531 = _T_2510 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294679.4]
  assign _T_2532 = _T_2530 | _T_2531; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294680.4]
  assign _T_2534 = _T_2532 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294682.4]
  assign _T_2535 = _T_2534 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294683.4]
  assign _T_2546 = _T_1057 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294700.4]
  assign _T_2547 = _T_1125 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294701.4]
  assign _T_2549 = _T_2547 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294703.4]
  assign _T_2551 = _T_2541 + _T_2546; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294705.4]
  assign _T_2552 = _T_2551 - _T_2549; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294706.4]
  assign _T_2553 = $unsigned(_T_2552); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294707.4]
  assign _T_2554 = _T_2553[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294708.4]
  assign _T_2555 = _T_2549 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294710.4]
  assign _T_2557 = _T_2555 | _T_2541; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294712.4]
  assign _T_2559 = _T_2557 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294714.4]
  assign _T_2560 = _T_2559 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294715.4]
  assign _T_2561 = _T_2546 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294720.4]
  assign _T_2562 = _T_2541 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294721.4]
  assign _T_2563 = _T_2561 | _T_2562; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294722.4]
  assign _T_2565 = _T_2563 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294724.4]
  assign _T_2566 = _T_2565 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294725.4]
  assign _T_2577 = _T_1058 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294742.4]
  assign _T_2578 = _T_1126 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294743.4]
  assign _T_2580 = _T_2578 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294745.4]
  assign _T_2582 = _T_2572 + _T_2577; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294747.4]
  assign _T_2583 = _T_2582 - _T_2580; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294748.4]
  assign _T_2584 = $unsigned(_T_2583); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294749.4]
  assign _T_2585 = _T_2584[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294750.4]
  assign _T_2586 = _T_2580 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294752.4]
  assign _T_2588 = _T_2586 | _T_2572; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294754.4]
  assign _T_2590 = _T_2588 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294756.4]
  assign _T_2591 = _T_2590 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294757.4]
  assign _T_2592 = _T_2577 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294762.4]
  assign _T_2593 = _T_2572 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294763.4]
  assign _T_2594 = _T_2592 | _T_2593; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294764.4]
  assign _T_2596 = _T_2594 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294766.4]
  assign _T_2597 = _T_2596 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294767.4]
  assign _T_2608 = _T_1059 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294784.4]
  assign _T_2609 = _T_1127 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294785.4]
  assign _T_2611 = _T_2609 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294787.4]
  assign _T_2613 = _T_2603 + _T_2608; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294789.4]
  assign _T_2614 = _T_2613 - _T_2611; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294790.4]
  assign _T_2615 = $unsigned(_T_2614); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294791.4]
  assign _T_2616 = _T_2615[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294792.4]
  assign _T_2617 = _T_2611 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294794.4]
  assign _T_2619 = _T_2617 | _T_2603; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294796.4]
  assign _T_2621 = _T_2619 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294798.4]
  assign _T_2622 = _T_2621 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294799.4]
  assign _T_2623 = _T_2608 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294804.4]
  assign _T_2624 = _T_2603 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294805.4]
  assign _T_2625 = _T_2623 | _T_2624; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294806.4]
  assign _T_2627 = _T_2625 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294808.4]
  assign _T_2628 = _T_2627 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294809.4]
  assign _T_2639 = _T_1060 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294826.4]
  assign _T_2640 = _T_1128 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294827.4]
  assign _T_2642 = _T_2640 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294829.4]
  assign _T_2644 = _T_2634 + _T_2639; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294831.4]
  assign _T_2645 = _T_2644 - _T_2642; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294832.4]
  assign _T_2646 = $unsigned(_T_2645); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294833.4]
  assign _T_2647 = _T_2646[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294834.4]
  assign _T_2648 = _T_2642 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294836.4]
  assign _T_2650 = _T_2648 | _T_2634; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294838.4]
  assign _T_2652 = _T_2650 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294840.4]
  assign _T_2653 = _T_2652 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294841.4]
  assign _T_2654 = _T_2639 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294846.4]
  assign _T_2655 = _T_2634 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294847.4]
  assign _T_2656 = _T_2654 | _T_2655; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294848.4]
  assign _T_2658 = _T_2656 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294850.4]
  assign _T_2659 = _T_2658 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294851.4]
  assign _T_2670 = _T_1061 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294868.4]
  assign _T_2671 = _T_1129 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294869.4]
  assign _T_2673 = _T_2671 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294871.4]
  assign _T_2675 = _T_2665 + _T_2670; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294873.4]
  assign _T_2676 = _T_2675 - _T_2673; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294874.4]
  assign _T_2677 = $unsigned(_T_2676); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294875.4]
  assign _T_2678 = _T_2677[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294876.4]
  assign _T_2679 = _T_2673 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294878.4]
  assign _T_2681 = _T_2679 | _T_2665; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294880.4]
  assign _T_2683 = _T_2681 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294882.4]
  assign _T_2684 = _T_2683 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294883.4]
  assign _T_2685 = _T_2670 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294888.4]
  assign _T_2686 = _T_2665 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294889.4]
  assign _T_2687 = _T_2685 | _T_2686; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294890.4]
  assign _T_2689 = _T_2687 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294892.4]
  assign _T_2690 = _T_2689 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294893.4]
  assign _T_2701 = _T_1062 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294910.4]
  assign _T_2702 = _T_1130 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294911.4]
  assign _T_2704 = _T_2702 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294913.4]
  assign _T_2706 = _T_2696 + _T_2701; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294915.4]
  assign _T_2707 = _T_2706 - _T_2704; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294916.4]
  assign _T_2708 = $unsigned(_T_2707); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294917.4]
  assign _T_2709 = _T_2708[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294918.4]
  assign _T_2710 = _T_2704 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294920.4]
  assign _T_2712 = _T_2710 | _T_2696; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294922.4]
  assign _T_2714 = _T_2712 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294924.4]
  assign _T_2715 = _T_2714 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294925.4]
  assign _T_2716 = _T_2701 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294930.4]
  assign _T_2717 = _T_2696 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294931.4]
  assign _T_2718 = _T_2716 | _T_2717; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294932.4]
  assign _T_2720 = _T_2718 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294934.4]
  assign _T_2721 = _T_2720 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294935.4]
  assign _T_2732 = _T_1063 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294952.4]
  assign _T_2733 = _T_1131 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294953.4]
  assign _T_2735 = _T_2733 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294955.4]
  assign _T_2737 = _T_2727 + _T_2732; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294957.4]
  assign _T_2738 = _T_2737 - _T_2735; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294958.4]
  assign _T_2739 = $unsigned(_T_2738); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294959.4]
  assign _T_2740 = _T_2739[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294960.4]
  assign _T_2741 = _T_2735 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294962.4]
  assign _T_2743 = _T_2741 | _T_2727; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294964.4]
  assign _T_2745 = _T_2743 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294966.4]
  assign _T_2746 = _T_2745 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294967.4]
  assign _T_2747 = _T_2732 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294972.4]
  assign _T_2748 = _T_2727 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294973.4]
  assign _T_2749 = _T_2747 | _T_2748; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294974.4]
  assign _T_2751 = _T_2749 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294976.4]
  assign _T_2752 = _T_2751 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294977.4]
  assign _T_2763 = _T_1064 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294994.4]
  assign _T_2764 = _T_1132 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294995.4]
  assign _T_2766 = _T_2764 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294997.4]
  assign _T_2768 = _T_2758 + _T_2763; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294999.4]
  assign _T_2769 = _T_2768 - _T_2766; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295000.4]
  assign _T_2770 = $unsigned(_T_2769); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295001.4]
  assign _T_2771 = _T_2770[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295002.4]
  assign _T_2772 = _T_2766 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295004.4]
  assign _T_2774 = _T_2772 | _T_2758; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295006.4]
  assign _T_2776 = _T_2774 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295008.4]
  assign _T_2777 = _T_2776 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295009.4]
  assign _T_2778 = _T_2763 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295014.4]
  assign _T_2779 = _T_2758 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295015.4]
  assign _T_2780 = _T_2778 | _T_2779; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295016.4]
  assign _T_2782 = _T_2780 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295018.4]
  assign _T_2783 = _T_2782 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295019.4]
  assign _T_2794 = _T_1065 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295036.4]
  assign _T_2795 = _T_1133 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295037.4]
  assign _T_2797 = _T_2795 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295039.4]
  assign _T_2799 = _T_2789 + _T_2794; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295041.4]
  assign _T_2800 = _T_2799 - _T_2797; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295042.4]
  assign _T_2801 = $unsigned(_T_2800); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295043.4]
  assign _T_2802 = _T_2801[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295044.4]
  assign _T_2803 = _T_2797 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295046.4]
  assign _T_2805 = _T_2803 | _T_2789; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295048.4]
  assign _T_2807 = _T_2805 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295050.4]
  assign _T_2808 = _T_2807 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295051.4]
  assign _T_2809 = _T_2794 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295056.4]
  assign _T_2810 = _T_2789 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295057.4]
  assign _T_2811 = _T_2809 | _T_2810; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295058.4]
  assign _T_2813 = _T_2811 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295060.4]
  assign _T_2814 = _T_2813 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295061.4]
  assign _T_2825 = _T_1066 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295078.4]
  assign _T_2826 = _T_1134 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295079.4]
  assign _T_2828 = _T_2826 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295081.4]
  assign _T_2830 = _T_2820 + _T_2825; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295083.4]
  assign _T_2831 = _T_2830 - _T_2828; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295084.4]
  assign _T_2832 = $unsigned(_T_2831); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295085.4]
  assign _T_2833 = _T_2832[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295086.4]
  assign _T_2834 = _T_2828 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295088.4]
  assign _T_2836 = _T_2834 | _T_2820; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295090.4]
  assign _T_2838 = _T_2836 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295092.4]
  assign _T_2839 = _T_2838 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295093.4]
  assign _T_2840 = _T_2825 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295098.4]
  assign _T_2841 = _T_2820 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295099.4]
  assign _T_2842 = _T_2840 | _T_2841; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295100.4]
  assign _T_2844 = _T_2842 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295102.4]
  assign _T_2845 = _T_2844 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295103.4]
  assign _T_2856 = _T_1067 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295120.4]
  assign _T_2857 = _T_1135 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295121.4]
  assign _T_2859 = _T_2857 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295123.4]
  assign _T_2861 = _T_2851 + _T_2856; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295125.4]
  assign _T_2862 = _T_2861 - _T_2859; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295126.4]
  assign _T_2863 = $unsigned(_T_2862); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295127.4]
  assign _T_2864 = _T_2863[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295128.4]
  assign _T_2865 = _T_2859 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295130.4]
  assign _T_2867 = _T_2865 | _T_2851; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295132.4]
  assign _T_2869 = _T_2867 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295134.4]
  assign _T_2870 = _T_2869 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295135.4]
  assign _T_2871 = _T_2856 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295140.4]
  assign _T_2872 = _T_2851 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295141.4]
  assign _T_2873 = _T_2871 | _T_2872; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295142.4]
  assign _T_2875 = _T_2873 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295144.4]
  assign _T_2876 = _T_2875 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295145.4]
  assign _T_2887 = _T_1068 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295162.4]
  assign _T_2888 = _T_1136 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295163.4]
  assign _T_2890 = _T_2888 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295165.4]
  assign _T_2892 = _T_2882 + _T_2887; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295167.4]
  assign _T_2893 = _T_2892 - _T_2890; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295168.4]
  assign _T_2894 = $unsigned(_T_2893); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295169.4]
  assign _T_2895 = _T_2894[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295170.4]
  assign _T_2896 = _T_2890 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295172.4]
  assign _T_2898 = _T_2896 | _T_2882; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295174.4]
  assign _T_2900 = _T_2898 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295176.4]
  assign _T_2901 = _T_2900 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295177.4]
  assign _T_2902 = _T_2887 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295182.4]
  assign _T_2903 = _T_2882 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295183.4]
  assign _T_2904 = _T_2902 | _T_2903; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295184.4]
  assign _T_2906 = _T_2904 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295186.4]
  assign _T_2907 = _T_2906 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295187.4]
  assign _T_2918 = _T_1069 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295204.4]
  assign _T_2919 = _T_1137 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295205.4]
  assign _T_2921 = _T_2919 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295207.4]
  assign _T_2923 = _T_2913 + _T_2918; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295209.4]
  assign _T_2924 = _T_2923 - _T_2921; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295210.4]
  assign _T_2925 = $unsigned(_T_2924); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295211.4]
  assign _T_2926 = _T_2925[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295212.4]
  assign _T_2927 = _T_2921 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295214.4]
  assign _T_2929 = _T_2927 | _T_2913; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295216.4]
  assign _T_2931 = _T_2929 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295218.4]
  assign _T_2932 = _T_2931 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295219.4]
  assign _T_2933 = _T_2918 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295224.4]
  assign _T_2934 = _T_2913 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295225.4]
  assign _T_2935 = _T_2933 | _T_2934; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295226.4]
  assign _T_2937 = _T_2935 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295228.4]
  assign _T_2938 = _T_2937 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295229.4]
  assign _T_2949 = _T_1070 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295246.4]
  assign _T_2950 = _T_1138 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295247.4]
  assign _T_2952 = _T_2950 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295249.4]
  assign _T_2954 = _T_2944 + _T_2949; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295251.4]
  assign _T_2955 = _T_2954 - _T_2952; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295252.4]
  assign _T_2956 = $unsigned(_T_2955); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295253.4]
  assign _T_2957 = _T_2956[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295254.4]
  assign _T_2958 = _T_2952 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295256.4]
  assign _T_2960 = _T_2958 | _T_2944; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295258.4]
  assign _T_2962 = _T_2960 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295260.4]
  assign _T_2963 = _T_2962 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295261.4]
  assign _T_2964 = _T_2949 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295266.4]
  assign _T_2965 = _T_2944 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295267.4]
  assign _T_2966 = _T_2964 | _T_2965; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295268.4]
  assign _T_2968 = _T_2966 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295270.4]
  assign _T_2969 = _T_2968 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295271.4]
  assign _T_2980 = _T_1071 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295288.4]
  assign _T_2981 = _T_1139 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295289.4]
  assign _T_2983 = _T_2981 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295291.4]
  assign _T_2985 = _T_2975 + _T_2980; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295293.4]
  assign _T_2986 = _T_2985 - _T_2983; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295294.4]
  assign _T_2987 = $unsigned(_T_2986); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295295.4]
  assign _T_2988 = _T_2987[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295296.4]
  assign _T_2989 = _T_2983 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295298.4]
  assign _T_2991 = _T_2989 | _T_2975; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295300.4]
  assign _T_2993 = _T_2991 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295302.4]
  assign _T_2994 = _T_2993 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295303.4]
  assign _T_2995 = _T_2980 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295308.4]
  assign _T_2996 = _T_2975 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295309.4]
  assign _T_2997 = _T_2995 | _T_2996; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295310.4]
  assign _T_2999 = _T_2997 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295312.4]
  assign _T_3000 = _T_2999 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295313.4]
  assign _T_3011 = _T_1072 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295330.4]
  assign _T_3012 = _T_1140 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295331.4]
  assign _T_3014 = _T_3012 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295333.4]
  assign _T_3016 = _T_3006 + _T_3011; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295335.4]
  assign _T_3017 = _T_3016 - _T_3014; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295336.4]
  assign _T_3018 = $unsigned(_T_3017); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295337.4]
  assign _T_3019 = _T_3018[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295338.4]
  assign _T_3020 = _T_3014 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295340.4]
  assign _T_3022 = _T_3020 | _T_3006; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295342.4]
  assign _T_3024 = _T_3022 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295344.4]
  assign _T_3025 = _T_3024 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295345.4]
  assign _T_3026 = _T_3011 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295350.4]
  assign _T_3027 = _T_3006 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295351.4]
  assign _T_3028 = _T_3026 | _T_3027; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295352.4]
  assign _T_3030 = _T_3028 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295354.4]
  assign _T_3031 = _T_3030 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295355.4]
  assign _T_3042 = _T_1073 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295372.4]
  assign _T_3043 = _T_1141 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295373.4]
  assign _T_3045 = _T_3043 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295375.4]
  assign _T_3047 = _T_3037 + _T_3042; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295377.4]
  assign _T_3048 = _T_3047 - _T_3045; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295378.4]
  assign _T_3049 = $unsigned(_T_3048); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295379.4]
  assign _T_3050 = _T_3049[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295380.4]
  assign _T_3051 = _T_3045 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295382.4]
  assign _T_3053 = _T_3051 | _T_3037; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295384.4]
  assign _T_3055 = _T_3053 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295386.4]
  assign _T_3056 = _T_3055 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295387.4]
  assign _T_3057 = _T_3042 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295392.4]
  assign _T_3058 = _T_3037 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295393.4]
  assign _T_3059 = _T_3057 | _T_3058; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295394.4]
  assign _T_3061 = _T_3059 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295396.4]
  assign _T_3062 = _T_3061 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295397.4]
  assign _T_3073 = _T_1074 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295414.4]
  assign _T_3074 = _T_1142 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295415.4]
  assign _T_3076 = _T_3074 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295417.4]
  assign _T_3078 = _T_3068 + _T_3073; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295419.4]
  assign _T_3079 = _T_3078 - _T_3076; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295420.4]
  assign _T_3080 = $unsigned(_T_3079); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295421.4]
  assign _T_3081 = _T_3080[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295422.4]
  assign _T_3082 = _T_3076 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295424.4]
  assign _T_3084 = _T_3082 | _T_3068; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295426.4]
  assign _T_3086 = _T_3084 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295428.4]
  assign _T_3087 = _T_3086 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295429.4]
  assign _T_3088 = _T_3073 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295434.4]
  assign _T_3089 = _T_3068 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295435.4]
  assign _T_3090 = _T_3088 | _T_3089; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295436.4]
  assign _T_3092 = _T_3090 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295438.4]
  assign _T_3093 = _T_3092 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295439.4]
  assign _T_3104 = _T_1075 & _T_1150; // @[ToAXI4.scala 229:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295456.4]
  assign _T_3105 = _T_1143 & _T_1144; // @[ToAXI4.scala 230:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295457.4]
  assign _T_3107 = _T_3105 & _T_1153; // @[ToAXI4.scala 230:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295459.4]
  assign _T_3109 = _T_3099 + _T_3104; // @[ToAXI4.scala 231:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295461.4]
  assign _T_3110 = _T_3109 - _T_3107; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295462.4]
  assign _T_3111 = $unsigned(_T_3110); // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295463.4]
  assign _T_3112 = _T_3111[0:0]; // @[ToAXI4.scala 231:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295464.4]
  assign _T_3113 = _T_3107 == 1'h0; // @[ToAXI4.scala 233:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295466.4]
  assign _T_3115 = _T_3113 | _T_3099; // @[ToAXI4.scala 233:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295468.4]
  assign _T_3117 = _T_3115 | reset; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295470.4]
  assign _T_3118 = _T_3117 == 1'h0; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295471.4]
  assign _T_3119 = _T_3104 == 1'h0; // @[ToAXI4.scala 234:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295476.4]
  assign _T_3120 = _T_3099 != 1'h1; // @[ToAXI4.scala 234:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295477.4]
  assign _T_3121 = _T_3119 | _T_3120; // @[ToAXI4.scala 234:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295478.4]
  assign _T_3123 = _T_3121 | reset; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295480.4]
  assign _T_3124 = _T_3123 == 1'h0; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295481.4]
  assign auto_in_a_ready = _T_970 & _T_973; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292136.4]
  assign auto_in_d_valid = _T_990 ? auto_out_r_valid : auto_out_b_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292136.4]
  assign auto_in_d_bits_opcode = _T_990 ? 3'h1 : 3'h0; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292136.4]
  assign auto_in_d_bits_size = _T_990 ? _T_923 : _T_925; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292136.4]
  assign auto_in_d_bits_source = _T_990 ? _T_922 : _T_924; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292136.4]
  assign auto_in_d_bits_denied = _T_990 ? _GEN_260 : _T_1002; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292136.4]
  assign auto_in_d_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292136.4]
  assign auto_in_d_bits_corrupt = _T_990 ? _T_1003 : 1'h0; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292136.4]
  assign auto_out_aw_valid = _T_948_valid & _T_948_bits_wen; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_id = Queue_1_io_deq_bits_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_addr = Queue_1_io_deq_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_len = Queue_1_io_deq_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_size = Queue_1_io_deq_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_burst = Queue_1_io_deq_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_lock = Queue_1_io_deq_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_cache = Queue_1_io_deq_bits_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_prot = Queue_1_io_deq_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_qos = Queue_1_io_deq_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_aw_bits_user = Queue_1_io_deq_bits_user; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_w_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_w_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_w_bits_strb = Queue_io_deq_bits_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_w_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_b_ready = auto_in_d_ready & _T_991; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_valid = _T_948_valid & _T_952; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_id = Queue_1_io_deq_bits_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_addr = Queue_1_io_deq_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_len = Queue_1_io_deq_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_size = Queue_1_io_deq_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_burst = Queue_1_io_deq_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_lock = Queue_1_io_deq_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_cache = Queue_1_io_deq_bits_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_prot = Queue_1_io_deq_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_qos = Queue_1_io_deq_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_ar_bits_user = Queue_1_io_deq_bits_user; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign auto_out_r_ready = auto_in_d_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292135.4]
  assign Queue_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292520.4]
  assign Queue_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292521.4]
  assign Queue_io_enq_valid = _T_983 & _T_971; // @[Decoupled.scala 294:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292522.4]
  assign Queue_io_enq_bits_data = auto_in_a_bits_data; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292525.4]
  assign Queue_io_enq_bits_strb = auto_in_a_bits_mask; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292524.4]
  assign Queue_io_enq_bits_last = _T_904 | _T_905; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292523.4]
  assign Queue_io_deq_ready = auto_out_w_ready; // @[Decoupled.scala 317:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292532.4]
  assign Queue_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292535.4]
  assign Queue_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292536.4]
  assign Queue_1_io_enq_valid = _T_976 & _T_979; // @[Decoupled.scala 294:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292537.4]
  assign Queue_1_io_enq_bits_id = 7'h7f == auto_in_a_bits_source ? 6'h3f : _GEN_128; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292548.4]
  assign Queue_1_io_enq_bits_addr = auto_in_a_bits_address; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292547.4]
  assign Queue_1_io_enq_bits_len = _T_964[10:3]; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292546.4]
  assign Queue_1_io_enq_bits_size = _T_966 ? 3'h3 : auto_in_a_bits_size; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292545.4]
  assign Queue_1_io_enq_bits_user = {{1'd0}, _T_921}; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292539.4]
  assign Queue_1_io_enq_bits_wen = _T_887 == 1'h0; // @[Decoupled.scala 295:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292538.4]
  assign Queue_1_io_deq_ready = _T_948_bits_wen ? auto_out_aw_ready : auto_out_ar_ready; // @[Decoupled.scala 317:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292563.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3099 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_3068 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_3037 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3006 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2975 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2944 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2913 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2882 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2851 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2820 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2789 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2758 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2727 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2696 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2665 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2634 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2603 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2572 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2541 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_2510 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2479 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2448 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2417 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2386 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2355 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_2324 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_2293 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_2262 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_2231 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_2200 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_2169 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_2138 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_2107 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_2076 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_2045 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_2014 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_1983 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_1952 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_1921 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_1890 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1859 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_1828 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_1797 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_1766 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_1735 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_1704 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_1673 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_1642 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1611 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_1580 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_1549 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1518 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1487 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_1456 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_1425 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1394 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_1363 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_1332 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_1301 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_1270 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_1239 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_1208 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_1177 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_1146 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_899 = _RAND_64[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_957 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_987 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_995 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_999 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_3099 <= 1'h0;
    end else begin
      _T_3099 <= _T_3112;
    end
    if (reset) begin
      _T_3068 <= 1'h0;
    end else begin
      _T_3068 <= _T_3081;
    end
    if (reset) begin
      _T_3037 <= 1'h0;
    end else begin
      _T_3037 <= _T_3050;
    end
    if (reset) begin
      _T_3006 <= 1'h0;
    end else begin
      _T_3006 <= _T_3019;
    end
    if (reset) begin
      _T_2975 <= 1'h0;
    end else begin
      _T_2975 <= _T_2988;
    end
    if (reset) begin
      _T_2944 <= 1'h0;
    end else begin
      _T_2944 <= _T_2957;
    end
    if (reset) begin
      _T_2913 <= 1'h0;
    end else begin
      _T_2913 <= _T_2926;
    end
    if (reset) begin
      _T_2882 <= 1'h0;
    end else begin
      _T_2882 <= _T_2895;
    end
    if (reset) begin
      _T_2851 <= 1'h0;
    end else begin
      _T_2851 <= _T_2864;
    end
    if (reset) begin
      _T_2820 <= 1'h0;
    end else begin
      _T_2820 <= _T_2833;
    end
    if (reset) begin
      _T_2789 <= 1'h0;
    end else begin
      _T_2789 <= _T_2802;
    end
    if (reset) begin
      _T_2758 <= 1'h0;
    end else begin
      _T_2758 <= _T_2771;
    end
    if (reset) begin
      _T_2727 <= 1'h0;
    end else begin
      _T_2727 <= _T_2740;
    end
    if (reset) begin
      _T_2696 <= 1'h0;
    end else begin
      _T_2696 <= _T_2709;
    end
    if (reset) begin
      _T_2665 <= 1'h0;
    end else begin
      _T_2665 <= _T_2678;
    end
    if (reset) begin
      _T_2634 <= 1'h0;
    end else begin
      _T_2634 <= _T_2647;
    end
    if (reset) begin
      _T_2603 <= 1'h0;
    end else begin
      _T_2603 <= _T_2616;
    end
    if (reset) begin
      _T_2572 <= 1'h0;
    end else begin
      _T_2572 <= _T_2585;
    end
    if (reset) begin
      _T_2541 <= 1'h0;
    end else begin
      _T_2541 <= _T_2554;
    end
    if (reset) begin
      _T_2510 <= 1'h0;
    end else begin
      _T_2510 <= _T_2523;
    end
    if (reset) begin
      _T_2479 <= 1'h0;
    end else begin
      _T_2479 <= _T_2492;
    end
    if (reset) begin
      _T_2448 <= 1'h0;
    end else begin
      _T_2448 <= _T_2461;
    end
    if (reset) begin
      _T_2417 <= 1'h0;
    end else begin
      _T_2417 <= _T_2430;
    end
    if (reset) begin
      _T_2386 <= 1'h0;
    end else begin
      _T_2386 <= _T_2399;
    end
    if (reset) begin
      _T_2355 <= 1'h0;
    end else begin
      _T_2355 <= _T_2368;
    end
    if (reset) begin
      _T_2324 <= 1'h0;
    end else begin
      _T_2324 <= _T_2337;
    end
    if (reset) begin
      _T_2293 <= 1'h0;
    end else begin
      _T_2293 <= _T_2306;
    end
    if (reset) begin
      _T_2262 <= 1'h0;
    end else begin
      _T_2262 <= _T_2275;
    end
    if (reset) begin
      _T_2231 <= 1'h0;
    end else begin
      _T_2231 <= _T_2244;
    end
    if (reset) begin
      _T_2200 <= 1'h0;
    end else begin
      _T_2200 <= _T_2213;
    end
    if (reset) begin
      _T_2169 <= 1'h0;
    end else begin
      _T_2169 <= _T_2182;
    end
    if (reset) begin
      _T_2138 <= 1'h0;
    end else begin
      _T_2138 <= _T_2151;
    end
    if (reset) begin
      _T_2107 <= 1'h0;
    end else begin
      _T_2107 <= _T_2120;
    end
    if (reset) begin
      _T_2076 <= 1'h0;
    end else begin
      _T_2076 <= _T_2089;
    end
    if (reset) begin
      _T_2045 <= 1'h0;
    end else begin
      _T_2045 <= _T_2058;
    end
    if (reset) begin
      _T_2014 <= 1'h0;
    end else begin
      _T_2014 <= _T_2027;
    end
    if (reset) begin
      _T_1983 <= 1'h0;
    end else begin
      _T_1983 <= _T_1996;
    end
    if (reset) begin
      _T_1952 <= 1'h0;
    end else begin
      _T_1952 <= _T_1965;
    end
    if (reset) begin
      _T_1921 <= 1'h0;
    end else begin
      _T_1921 <= _T_1934;
    end
    if (reset) begin
      _T_1890 <= 1'h0;
    end else begin
      _T_1890 <= _T_1903;
    end
    if (reset) begin
      _T_1859 <= 1'h0;
    end else begin
      _T_1859 <= _T_1872;
    end
    if (reset) begin
      _T_1828 <= 1'h0;
    end else begin
      _T_1828 <= _T_1841;
    end
    if (reset) begin
      _T_1797 <= 1'h0;
    end else begin
      _T_1797 <= _T_1810;
    end
    if (reset) begin
      _T_1766 <= 1'h0;
    end else begin
      _T_1766 <= _T_1779;
    end
    if (reset) begin
      _T_1735 <= 1'h0;
    end else begin
      _T_1735 <= _T_1748;
    end
    if (reset) begin
      _T_1704 <= 1'h0;
    end else begin
      _T_1704 <= _T_1717;
    end
    if (reset) begin
      _T_1673 <= 1'h0;
    end else begin
      _T_1673 <= _T_1686;
    end
    if (reset) begin
      _T_1642 <= 1'h0;
    end else begin
      _T_1642 <= _T_1655;
    end
    if (reset) begin
      _T_1611 <= 1'h0;
    end else begin
      _T_1611 <= _T_1624;
    end
    if (reset) begin
      _T_1580 <= 1'h0;
    end else begin
      _T_1580 <= _T_1593;
    end
    if (reset) begin
      _T_1549 <= 1'h0;
    end else begin
      _T_1549 <= _T_1562;
    end
    if (reset) begin
      _T_1518 <= 1'h0;
    end else begin
      _T_1518 <= _T_1531;
    end
    if (reset) begin
      _T_1487 <= 1'h0;
    end else begin
      _T_1487 <= _T_1500;
    end
    if (reset) begin
      _T_1456 <= 1'h0;
    end else begin
      _T_1456 <= _T_1469;
    end
    if (reset) begin
      _T_1425 <= 1'h0;
    end else begin
      _T_1425 <= _T_1438;
    end
    if (reset) begin
      _T_1394 <= 1'h0;
    end else begin
      _T_1394 <= _T_1407;
    end
    if (reset) begin
      _T_1363 <= 1'h0;
    end else begin
      _T_1363 <= _T_1376;
    end
    if (reset) begin
      _T_1332 <= 1'h0;
    end else begin
      _T_1332 <= _T_1345;
    end
    if (reset) begin
      _T_1301 <= 1'h0;
    end else begin
      _T_1301 <= _T_1314;
    end
    if (reset) begin
      _T_1270 <= 1'h0;
    end else begin
      _T_1270 <= _T_1283;
    end
    if (reset) begin
      _T_1239 <= 1'h0;
    end else begin
      _T_1239 <= _T_1252;
    end
    if (reset) begin
      _T_1208 <= 1'h0;
    end else begin
      _T_1208 <= _T_1221;
    end
    if (reset) begin
      _T_1177 <= 1'h0;
    end else begin
      _T_1177 <= _T_1190;
    end
    if (reset) begin
      _T_1146 <= 1'h0;
    end else begin
      _T_1146 <= _T_1159;
    end
    if (reset) begin
      _T_899 <= 4'h0;
    end else begin
      if (_T_889) begin
        if (_T_903) begin
          if (_T_888) begin
            _T_899 <= _T_894;
          end else begin
            _T_899 <= 4'h0;
          end
        end else begin
          _T_899 <= _T_902;
        end
      end
    end
    if (reset) begin
      _T_957 <= 1'h0;
    end else begin
      if (_T_889) begin
        _T_957 <= _T_959;
      end
    end
    if (reset) begin
      _T_987 <= 1'h0;
    end else begin
      if (_T_988) begin
        _T_987 <= _T_989;
      end
    end
    if (reset) begin
      _T_995 <= 1'h1;
    end else begin
      if (_T_988) begin
        _T_995 <= auto_out_r_bits_last;
      end
    end
    if (_T_995) begin
      _T_999 <= _T_997;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:125 assert (a_source  < UInt(BigInt(1) << sourceBits))\n"); // @[ToAXI4.scala 125:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292497.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[ToAXI4.scala 125:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292498.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:126 assert (a_size    < UInt(BigInt(1) << sizeBits))\n"); // @[ToAXI4.scala 126:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292505.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[ToAXI4.scala 126:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292506.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1165) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292827.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1165) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292828.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1171) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292837.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1171) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292838.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1196) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292869.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1196) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292870.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1202) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292879.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1202) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292880.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1227) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292911.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1227) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292912.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1233) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292921.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1233) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292922.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1258) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292953.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1258) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292954.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1264) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292963.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1264) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292964.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1289) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292995.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1289) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@292996.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1295) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293005.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1295) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293006.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1320) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293037.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1320) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293038.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1326) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293047.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1326) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293048.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1351) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293079.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1351) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293080.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1357) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293089.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1357) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293090.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1382) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293121.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1382) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293122.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1388) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293131.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1388) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293132.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1413) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293163.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1413) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293164.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1419) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293173.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1419) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293174.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1444) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293205.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1444) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293206.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1450) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293215.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1450) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293216.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1475) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293247.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1475) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293248.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1481) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293257.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1481) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293258.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1506) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293289.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1506) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293290.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1512) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293299.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1512) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293300.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1537) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293331.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1537) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293332.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1543) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293341.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1543) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293342.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1568) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293373.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1568) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293374.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1574) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293383.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1574) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293384.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1599) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293415.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1599) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293416.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293425.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293426.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1630) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293457.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1630) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293458.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1636) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293467.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1636) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293468.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1661) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293499.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1661) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293500.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1667) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293509.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1667) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293510.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1692) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293541.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1692) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293542.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1698) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293551.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1698) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293552.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1723) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293583.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1723) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293584.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1729) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293593.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1729) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293594.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1754) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293625.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1754) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293626.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1760) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293635.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1760) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293636.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1785) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293667.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1785) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293668.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1791) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293677.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1791) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293678.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1816) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293709.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1816) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293710.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1822) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293719.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1822) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293720.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1847) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293751.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1847) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293752.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1853) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293761.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1853) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293762.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1878) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293793.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1878) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293794.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1884) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293803.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1884) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293804.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1909) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293835.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1909) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293836.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1915) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293845.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1915) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293846.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1940) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293877.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1940) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293878.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1946) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293887.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1946) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293888.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1971) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293919.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1971) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293920.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1977) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293929.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1977) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293930.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2002) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293961.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2002) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293962.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2008) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293971.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2008) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@293972.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2033) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294003.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2033) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294004.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2039) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294013.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2039) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294014.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2064) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294045.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2064) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294046.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2070) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294055.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2070) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294056.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2095) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294087.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2095) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294088.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2101) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294097.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2101) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294098.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2126) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294129.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2126) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294130.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2132) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294139.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2132) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294140.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2157) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294171.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2157) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294172.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2163) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294181.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2163) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294182.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294213.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294214.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2194) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294223.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2194) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294224.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2219) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294255.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2219) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294256.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2225) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294265.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2225) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294266.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2250) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294297.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2250) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294298.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2256) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294307.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2256) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294308.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2281) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294339.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2281) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294340.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2287) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294349.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2287) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294350.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2312) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294381.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2312) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294382.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2318) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294391.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2318) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294392.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2343) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294423.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2343) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294424.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2349) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294433.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2349) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294434.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2374) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294465.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2374) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294466.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2380) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294475.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2380) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294476.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2405) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294507.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2405) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294508.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2411) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294517.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2411) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294518.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2436) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294549.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2436) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294550.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2442) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294559.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2442) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294560.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2467) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294591.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2467) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294592.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2473) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294601.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2473) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294602.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2498) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294633.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2498) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294634.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2504) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294643.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2504) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294644.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2529) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294675.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2529) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294676.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2535) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294685.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2535) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294686.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2560) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294717.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2560) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294718.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2566) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294727.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2566) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294728.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2591) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294759.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2591) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294760.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2597) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294769.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2597) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294770.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2622) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294801.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2622) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294802.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2628) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294811.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2628) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294812.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2653) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294843.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2653) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294844.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2659) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294853.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2659) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294854.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2684) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294885.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2684) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294886.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2690) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294895.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2690) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294896.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2715) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294927.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2715) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294928.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2721) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294937.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2721) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294938.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2746) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294969.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2746) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294970.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2752) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294979.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2752) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@294980.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2777) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295011.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2777) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295012.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2783) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295021.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2783) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295022.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2808) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295053.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2808) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295054.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295063.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295064.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2839) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295095.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2839) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295096.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2845) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295105.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2845) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295106.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2870) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295137.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2870) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295138.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2876) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295147.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2876) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295148.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295179.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295180.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2907) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295189.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2907) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295190.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2932) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295221.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2932) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295222.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2938) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295231.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2938) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295232.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2963) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295263.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2963) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295264.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2969) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295273.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2969) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295274.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2994) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295305.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2994) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295306.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3000) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295315.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3000) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295316.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3025) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295347.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3025) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295348.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3031) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295357.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3031) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295358.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3056) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295389.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3056) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295390.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3062) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295399.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3062) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295400.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3087) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295431.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3087) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295432.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3093) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295441.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3093) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295442.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3118) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295473.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3118) begin
          $fatal; // @[ToAXI4.scala 233:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295474.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3124) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295483.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3124) begin
          $fatal; // @[ToAXI4.scala 234:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295484.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295498.2]
  output        auto_in_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_in_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [5:0]  auto_in_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [31:0] auto_in_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_in_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [10:0] auto_in_aw_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_in_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_in_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [63:0] auto_in_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [7:0]  auto_in_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_in_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_in_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_in_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [5:0]  auto_in_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [1:0]  auto_in_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [10:0] auto_in_b_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_in_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_in_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [5:0]  auto_in_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [31:0] auto_in_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_in_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [10:0] auto_in_ar_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_in_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_in_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [5:0]  auto_in_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [63:0] auto_in_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [1:0]  auto_in_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [10:0] auto_in_r_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_in_r_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_out_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_out_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [3:0]  auto_out_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [31:0] auto_out_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [7:0]  auto_out_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [2:0]  auto_out_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_out_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [12:0] auto_out_aw_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_out_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_out_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [63:0] auto_out_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [7:0]  auto_out_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_out_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_out_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_out_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [3:0]  auto_out_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [12:0] auto_out_b_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_out_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_out_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [3:0]  auto_out_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [31:0] auto_out_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [7:0]  auto_out_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [2:0]  auto_out_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_out_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output [12:0] auto_out_ar_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  output        auto_out_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_out_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [3:0]  auto_out_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [63:0] auto_out_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input  [12:0] auto_out_r_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
  input         auto_out_r_bits_last // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295501.4]
);
  wire [1:0] _T_221; // @[IdIndexer.scala 56:81:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295517.4]
  wire [1:0] _T_223; // @[IdIndexer.scala 57:81:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295520.4]
  wire [16:0] _T_227; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295527.4]
  wire [16:0] _T_228; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295529.4]
  assign _T_221 = auto_in_ar_bits_id[5:4]; // @[IdIndexer.scala 56:81:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295517.4]
  assign _T_223 = auto_in_aw_bits_id[5:4]; // @[IdIndexer.scala 57:81:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295520.4]
  assign _T_227 = {auto_out_r_bits_user,auto_out_r_bits_id}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295527.4]
  assign _T_228 = {auto_out_b_bits_user,auto_out_b_bits_id}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295529.4]
  assign auto_in_aw_ready = auto_out_aw_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_b_bits_id = _T_228[5:0]; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_b_bits_user = auto_out_b_bits_user[12:2]; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_r_bits_id = _T_227[5:0]; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_r_bits_user = auto_out_r_bits_user[12:2]; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295511.4]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id[3:0]; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_aw_bits_user = {auto_in_aw_bits_user,_T_223}; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id[3:0]; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_ar_bits_user = {auto_in_ar_bits_user,_T_221}; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295510.4]
endmodule
module Queue_46( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295532.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295533.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295534.4]
  output        io_enq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  input         io_enq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  input  [3:0]  io_enq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  input  [63:0] io_enq_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  input  [1:0]  io_enq_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  input  [12:0] io_enq_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  input         io_enq_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  input         io_deq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  output        io_deq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  output [3:0]  io_deq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  output [63:0] io_deq_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  output [1:0]  io_deq_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  output [12:0] io_deq_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
  output        io_deq_bits_last // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295535.4]
);
  reg [3:0] _T_35_id [0:7]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [31:0] _RAND_0;
  wire [3:0] _T_35_id__T_58_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_id__T_58_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [3:0] _T_35_id__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_id__T_50_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_id__T_50_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_id__T_50_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [63:0] _T_35_data [0:7]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [63:0] _RAND_1;
  wire [63:0] _T_35_data__T_58_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_data__T_58_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [63:0] _T_35_data__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_data__T_50_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_data__T_50_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_data__T_50_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [1:0] _T_35_resp [0:7]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [31:0] _RAND_2;
  wire [1:0] _T_35_resp__T_58_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_resp__T_58_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [1:0] _T_35_resp__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_resp__T_50_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_resp__T_50_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_resp__T_50_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [12:0] _T_35_user [0:7]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [31:0] _RAND_3;
  wire [12:0] _T_35_user__T_58_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_user__T_58_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [12:0] _T_35_user__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_user__T_50_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_user__T_50_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_user__T_50_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg  _T_35_last [0:7]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [31:0] _RAND_4;
  wire  _T_35_last__T_58_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_last__T_58_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_last__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire [2:0] _T_35_last__T_50_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_last__T_50_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  wire  _T_35_last__T_50_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  reg [2:0] value; // @[Counter.scala 26:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295541.4]
  reg [31:0] _RAND_5;
  reg [2:0] value_1; // @[Counter.scala 26:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295542.4]
  reg [31:0] _RAND_6;
  reg  _T_39; // @[Decoupled.scala 217:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295543.4]
  reg [31:0] _RAND_7;
  wire  _T_40; // @[Decoupled.scala 219:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295544.4]
  wire  _T_41; // @[Decoupled.scala 220:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295545.4]
  wire  _T_42; // @[Decoupled.scala 220:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295546.4]
  wire  _T_43; // @[Decoupled.scala 221:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295547.4]
  wire  _T_44; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295548.4]
  wire  _T_47; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295552.4]
  wire [2:0] _T_52; // @[Counter.scala 35:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295561.6]
  wire [2:0] _T_54; // @[Counter.scala 35:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295567.6]
  wire  _T_55; // @[Decoupled.scala 232:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295570.4]
  assign _T_35_id__T_58_addr = value_1;
  assign _T_35_id__T_58_data = _T_35_id[_T_35_id__T_58_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  assign _T_35_id__T_50_data = io_enq_bits_id;
  assign _T_35_id__T_50_addr = value;
  assign _T_35_id__T_50_mask = 1'h1;
  assign _T_35_id__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_data__T_58_addr = value_1;
  assign _T_35_data__T_58_data = _T_35_data[_T_35_data__T_58_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  assign _T_35_data__T_50_data = io_enq_bits_data;
  assign _T_35_data__T_50_addr = value;
  assign _T_35_data__T_50_mask = 1'h1;
  assign _T_35_data__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_resp__T_58_addr = value_1;
  assign _T_35_resp__T_58_data = _T_35_resp[_T_35_resp__T_58_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  assign _T_35_resp__T_50_data = io_enq_bits_resp;
  assign _T_35_resp__T_50_addr = value;
  assign _T_35_resp__T_50_mask = 1'h1;
  assign _T_35_resp__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_user__T_58_addr = value_1;
  assign _T_35_user__T_58_data = _T_35_user[_T_35_user__T_58_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  assign _T_35_user__T_50_data = io_enq_bits_user;
  assign _T_35_user__T_50_addr = value;
  assign _T_35_user__T_50_mask = 1'h1;
  assign _T_35_user__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_last__T_58_addr = value_1;
  assign _T_35_last__T_58_data = _T_35_last[_T_35_last__T_58_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
  assign _T_35_last__T_50_data = io_enq_bits_last;
  assign _T_35_last__T_50_addr = value;
  assign _T_35_last__T_50_mask = 1'h1;
  assign _T_35_last__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_40 = value == value_1; // @[Decoupled.scala 219:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295544.4]
  assign _T_41 = _T_39 == 1'h0; // @[Decoupled.scala 220:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295545.4]
  assign _T_42 = _T_40 & _T_41; // @[Decoupled.scala 220:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295546.4]
  assign _T_43 = _T_40 & _T_39; // @[Decoupled.scala 221:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295547.4]
  assign _T_44 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295548.4]
  assign _T_47 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295552.4]
  assign _T_52 = value + 3'h1; // @[Counter.scala 35:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295561.6]
  assign _T_54 = value_1 + 3'h1; // @[Counter.scala 35:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295567.6]
  assign _T_55 = _T_44 != _T_47; // @[Decoupled.scala 232:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295570.4]
  assign io_enq_ready = _T_43 == 1'h0; // @[Decoupled.scala 237:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295577.4]
  assign io_deq_valid = _T_42 == 1'h0; // @[Decoupled.scala 236:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295575.4]
  assign io_deq_bits_id = _T_35_id__T_58_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295579.4]
  assign io_deq_bits_data = _T_35_data__T_58_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295579.4]
  assign io_deq_bits_resp = _T_35_resp__T_58_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295579.4]
  assign io_deq_bits_user = _T_35_user__T_58_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295579.4]
  assign io_deq_bits_last = _T_35_last__T_58_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295579.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_35_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_35_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_35_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_35_user[initvar] = _RAND_3[12:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_35_last[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_1 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_39 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35_id__T_50_en & _T_35_id__T_50_mask) begin
      _T_35_id[_T_35_id__T_50_addr] <= _T_35_id__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
    end
    if(_T_35_data__T_50_en & _T_35_data__T_50_mask) begin
      _T_35_data[_T_35_data__T_50_addr] <= _T_35_data__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
    end
    if(_T_35_resp__T_50_en & _T_35_resp__T_50_mask) begin
      _T_35_resp[_T_35_resp__T_50_addr] <= _T_35_resp__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
    end
    if(_T_35_user__T_50_en & _T_35_user__T_50_mask) begin
      _T_35_user[_T_35_user__T_50_addr] <= _T_35_user__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
    end
    if(_T_35_last__T_50_en & _T_35_last__T_50_mask) begin
      _T_35_last[_T_35_last__T_50_addr] <= _T_35_last__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@295540.4]
    end
    if (reset) begin
      value <= 3'h0;
    end else begin
      if (_T_44) begin
        value <= _T_52;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (_T_47) begin
        value_1 <= _T_54;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_55) begin
        _T_39 <= _T_44;
      end
    end
  end
endmodule
module AXI4Deinterleaver( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296412.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296413.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296414.4]
  output        auto_in_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_in_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [3:0]  auto_in_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [31:0] auto_in_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_in_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [12:0] auto_in_aw_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_in_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_in_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [63:0] auto_in_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [7:0]  auto_in_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_in_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_in_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_in_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [3:0]  auto_in_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [1:0]  auto_in_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [12:0] auto_in_b_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_in_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_in_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [3:0]  auto_in_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [31:0] auto_in_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_in_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [12:0] auto_in_ar_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_in_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_in_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [3:0]  auto_in_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [63:0] auto_in_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [1:0]  auto_in_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [12:0] auto_in_r_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_in_r_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_out_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_out_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [3:0]  auto_out_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [31:0] auto_out_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [7:0]  auto_out_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [2:0]  auto_out_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_out_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [12:0] auto_out_aw_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_out_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_out_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [63:0] auto_out_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [7:0]  auto_out_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_out_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_out_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_out_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [3:0]  auto_out_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [12:0] auto_out_b_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_out_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_out_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [3:0]  auto_out_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [31:0] auto_out_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [7:0]  auto_out_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [2:0]  auto_out_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_out_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output [12:0] auto_out_ar_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  output        auto_out_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_out_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [3:0]  auto_out_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [63:0] auto_out_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input  [12:0] auto_out_r_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
  input         auto_out_r_bits_last // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296415.4]
);
  wire  Queue_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire  Queue_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire  Queue_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire  Queue_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire [3:0] Queue_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire [63:0] Queue_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire [1:0] Queue_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire [12:0] Queue_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire  Queue_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire  Queue_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire  Queue_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire [3:0] Queue_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire [63:0] Queue_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire [1:0] Queue_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire [12:0] Queue_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire  Queue_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
  wire  Queue_1_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire  Queue_1_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire  Queue_1_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire  Queue_1_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire [3:0] Queue_1_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire [63:0] Queue_1_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire [1:0] Queue_1_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire [12:0] Queue_1_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire  Queue_1_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire  Queue_1_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire  Queue_1_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire [3:0] Queue_1_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire [63:0] Queue_1_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire [1:0] Queue_1_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire [12:0] Queue_1_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire  Queue_1_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
  wire  Queue_2_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire  Queue_2_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire  Queue_2_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire  Queue_2_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire [3:0] Queue_2_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire [63:0] Queue_2_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire [1:0] Queue_2_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire [12:0] Queue_2_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire  Queue_2_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire  Queue_2_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire  Queue_2_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire [3:0] Queue_2_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire [63:0] Queue_2_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire [1:0] Queue_2_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire [12:0] Queue_2_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire  Queue_2_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
  wire  Queue_3_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire  Queue_3_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire  Queue_3_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire  Queue_3_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire [3:0] Queue_3_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire [63:0] Queue_3_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire [1:0] Queue_3_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire [12:0] Queue_3_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire  Queue_3_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire  Queue_3_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire  Queue_3_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire [3:0] Queue_3_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire [63:0] Queue_3_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire [1:0] Queue_3_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire [12:0] Queue_3_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire  Queue_3_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
  wire  Queue_4_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire  Queue_4_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire  Queue_4_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire  Queue_4_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire [3:0] Queue_4_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire [63:0] Queue_4_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire [1:0] Queue_4_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire [12:0] Queue_4_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire  Queue_4_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire  Queue_4_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire  Queue_4_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire [3:0] Queue_4_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire [63:0] Queue_4_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire [1:0] Queue_4_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire [12:0] Queue_4_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire  Queue_4_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
  wire  Queue_5_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire  Queue_5_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire  Queue_5_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire  Queue_5_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire [3:0] Queue_5_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire [63:0] Queue_5_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire [1:0] Queue_5_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire [12:0] Queue_5_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire  Queue_5_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire  Queue_5_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire  Queue_5_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire [3:0] Queue_5_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire [63:0] Queue_5_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire [1:0] Queue_5_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire [12:0] Queue_5_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire  Queue_5_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
  wire  Queue_6_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire  Queue_6_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire  Queue_6_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire  Queue_6_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire [3:0] Queue_6_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire [63:0] Queue_6_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire [1:0] Queue_6_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire [12:0] Queue_6_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire  Queue_6_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire  Queue_6_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire  Queue_6_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire [3:0] Queue_6_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire [63:0] Queue_6_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire [1:0] Queue_6_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire [12:0] Queue_6_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire  Queue_6_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
  wire  Queue_7_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire  Queue_7_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire  Queue_7_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire  Queue_7_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire [3:0] Queue_7_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire [63:0] Queue_7_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire [1:0] Queue_7_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire [12:0] Queue_7_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire  Queue_7_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire  Queue_7_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire  Queue_7_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire [3:0] Queue_7_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire [63:0] Queue_7_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire [1:0] Queue_7_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire [12:0] Queue_7_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire  Queue_7_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
  wire  Queue_8_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire  Queue_8_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire  Queue_8_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire  Queue_8_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire [3:0] Queue_8_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire [63:0] Queue_8_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire [1:0] Queue_8_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire [12:0] Queue_8_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire  Queue_8_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire  Queue_8_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire  Queue_8_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire [3:0] Queue_8_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire [63:0] Queue_8_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire [1:0] Queue_8_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire [12:0] Queue_8_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire  Queue_8_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
  wire  Queue_9_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire  Queue_9_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire  Queue_9_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire  Queue_9_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire [3:0] Queue_9_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire [63:0] Queue_9_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire [1:0] Queue_9_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire [12:0] Queue_9_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire  Queue_9_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire  Queue_9_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire  Queue_9_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire [3:0] Queue_9_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire [63:0] Queue_9_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire [1:0] Queue_9_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire [12:0] Queue_9_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire  Queue_9_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
  wire  Queue_10_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire  Queue_10_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire  Queue_10_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire  Queue_10_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire [3:0] Queue_10_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire [63:0] Queue_10_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire [1:0] Queue_10_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire [12:0] Queue_10_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire  Queue_10_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire  Queue_10_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire  Queue_10_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire [3:0] Queue_10_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire [63:0] Queue_10_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire [1:0] Queue_10_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire [12:0] Queue_10_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire  Queue_10_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
  wire  Queue_11_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire  Queue_11_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire  Queue_11_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire  Queue_11_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire [3:0] Queue_11_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire [63:0] Queue_11_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire [1:0] Queue_11_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire [12:0] Queue_11_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire  Queue_11_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire  Queue_11_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire  Queue_11_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire [3:0] Queue_11_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire [63:0] Queue_11_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire [1:0] Queue_11_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire [12:0] Queue_11_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire  Queue_11_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
  wire  Queue_12_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire  Queue_12_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire  Queue_12_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire  Queue_12_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire [3:0] Queue_12_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire [63:0] Queue_12_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire [1:0] Queue_12_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire [12:0] Queue_12_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire  Queue_12_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire  Queue_12_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire  Queue_12_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire [3:0] Queue_12_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire [63:0] Queue_12_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire [1:0] Queue_12_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire [12:0] Queue_12_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire  Queue_12_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
  wire  Queue_13_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire  Queue_13_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire  Queue_13_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire  Queue_13_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire [3:0] Queue_13_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire [63:0] Queue_13_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire [1:0] Queue_13_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire [12:0] Queue_13_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire  Queue_13_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire  Queue_13_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire  Queue_13_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire [3:0] Queue_13_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire [63:0] Queue_13_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire [1:0] Queue_13_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire [12:0] Queue_13_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire  Queue_13_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
  wire  Queue_14_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire  Queue_14_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire  Queue_14_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire  Queue_14_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire [3:0] Queue_14_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire [63:0] Queue_14_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire [1:0] Queue_14_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire [12:0] Queue_14_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire  Queue_14_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire  Queue_14_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire  Queue_14_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire [3:0] Queue_14_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire [63:0] Queue_14_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire [1:0] Queue_14_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire [12:0] Queue_14_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire  Queue_14_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
  wire  Queue_15_clock; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire  Queue_15_reset; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire  Queue_15_io_enq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire  Queue_15_io_enq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire [3:0] Queue_15_io_enq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire [63:0] Queue_15_io_enq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire [1:0] Queue_15_io_enq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire [12:0] Queue_15_io_enq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire  Queue_15_io_enq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire  Queue_15_io_deq_ready; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire  Queue_15_io_deq_valid; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire [3:0] Queue_15_io_deq_bits_id; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire [63:0] Queue_15_io_deq_bits_data; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire [1:0] Queue_15_io_deq_bits_resp; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire [12:0] Queue_15_io_deq_bits_user; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  wire  Queue_15_io_deq_bits_last; // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
  reg  _T_222; // @[Deinterleaver.scala 50:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296494.4]
  reg [31:0] _RAND_0;
  reg [3:0] _T_224; // @[Deinterleaver.scala 51:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296495.4]
  reg [31:0] _RAND_1;
  wire [15:0] _T_226; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296497.4]
  wire [15:0] _T_229; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296500.4]
  reg [3:0] _T_232; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296502.4]
  reg [31:0] _RAND_2;
  wire  _T_234; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296505.4]
  wire  _T_826_15; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297288.4]
  wire  _T_826_14; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297287.4]
  wire  _T_826_13; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297286.4]
  wire  _T_826_12; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297285.4]
  wire  _T_826_11; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297284.4]
  wire  _T_826_10; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297283.4]
  wire  _T_826_9; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297282.4]
  wire  _T_826_8; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297281.4]
  wire  _T_826_7; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297280.4]
  wire  _T_826_6; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297279.4]
  wire  _T_826_5; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297278.4]
  wire  _T_826_4; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297277.4]
  wire  _T_826_3; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297276.4]
  wire  _T_826_2; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297275.4]
  wire  _T_826_1; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297274.4]
  wire  _T_826_0; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297273.4]
  wire  _GEN_83; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_84; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_85; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_86; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_87; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_88; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_89; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_90; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_91; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_92; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_93; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_94; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_95; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_96; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _GEN_97; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  wire  _T_235; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296506.4]
  wire  _T_236; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296507.4]
  wire  _T_237; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296508.4]
  wire  _T_238; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296509.4]
  wire  _T_239; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296510.4]
  wire  _T_240; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296511.4]
  wire  _T_755_15_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  wire  _T_755_14_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  wire  _T_755_13_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  wire  _T_755_12_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  wire  _T_755_11_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  wire  _T_755_10_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  wire  _T_755_9_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  wire  _T_755_8_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  wire  _T_755_7_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  wire  _T_755_6_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  wire  _T_755_5_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  wire  _T_755_4_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  wire  _T_755_3_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  wire  _T_755_2_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  wire  _T_755_1_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  wire  _T_755_0_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  wire  _GEN_11; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_16; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_21; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_26; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_31; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_36; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_41; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_46; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_51; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_56; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_61; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_66; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_71; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_76; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _GEN_81; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire  _T_241; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296512.4]
  wire [3:0] _GEN_98; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296513.4]
  wire [3:0] _T_243; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296514.4]
  wire [3:0] _GEN_99; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296515.4]
  wire [4:0] _T_244; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296515.4]
  wire [4:0] _T_245; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296516.4]
  wire [3:0] _T_246; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296517.4]
  wire  _T_247; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296520.4]
  wire  _T_248; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296521.4]
  wire  _T_249; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296522.4]
  wire  _T_251; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296524.4]
  wire  _T_252; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296525.4]
  wire  _T_253; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296530.4]
  wire  _T_254; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296531.4]
  wire  _T_255; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296532.4]
  wire  _T_257; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296534.4]
  wire  _T_258; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296535.4]
  wire  _T_259; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296540.4]
  reg [3:0] _T_261; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296541.4]
  reg [31:0] _RAND_3;
  wire  _T_263; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296544.4]
  wire  _T_265; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296546.4]
  wire  _T_266; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296547.4]
  wire  _T_267; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296548.4]
  wire  _T_269; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296550.4]
  wire  _T_270; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296551.4]
  wire [3:0] _GEN_100; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296552.4]
  wire [3:0] _T_272; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296553.4]
  wire [3:0] _GEN_101; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296554.4]
  wire [4:0] _T_273; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296554.4]
  wire [4:0] _T_274; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296555.4]
  wire [3:0] _T_275; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296556.4]
  wire  _T_276; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296559.4]
  wire  _T_277; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296560.4]
  wire  _T_278; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296561.4]
  wire  _T_280; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296563.4]
  wire  _T_281; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296564.4]
  wire  _T_282; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296569.4]
  wire  _T_283; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296570.4]
  wire  _T_284; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296571.4]
  wire  _T_286; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296573.4]
  wire  _T_287; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296574.4]
  wire  _T_288; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296579.4]
  reg [3:0] _T_290; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296580.4]
  reg [31:0] _RAND_4;
  wire  _T_292; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296583.4]
  wire  _T_294; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296585.4]
  wire  _T_295; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296586.4]
  wire  _T_296; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296587.4]
  wire  _T_298; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296589.4]
  wire  _T_299; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296590.4]
  wire [3:0] _GEN_102; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296591.4]
  wire [3:0] _T_301; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296592.4]
  wire [3:0] _GEN_103; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296593.4]
  wire [4:0] _T_302; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296593.4]
  wire [4:0] _T_303; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296594.4]
  wire [3:0] _T_304; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296595.4]
  wire  _T_305; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296598.4]
  wire  _T_306; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296599.4]
  wire  _T_307; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296600.4]
  wire  _T_309; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296602.4]
  wire  _T_310; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296603.4]
  wire  _T_311; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296608.4]
  wire  _T_312; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296609.4]
  wire  _T_313; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296610.4]
  wire  _T_315; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296612.4]
  wire  _T_316; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296613.4]
  wire  _T_317; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296618.4]
  reg [3:0] _T_319; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296619.4]
  reg [31:0] _RAND_5;
  wire  _T_321; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296622.4]
  wire  _T_323; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296624.4]
  wire  _T_324; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296625.4]
  wire  _T_325; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296626.4]
  wire  _T_327; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296628.4]
  wire  _T_328; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296629.4]
  wire [3:0] _GEN_104; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296630.4]
  wire [3:0] _T_330; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296631.4]
  wire [3:0] _GEN_105; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296632.4]
  wire [4:0] _T_331; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296632.4]
  wire [4:0] _T_332; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296633.4]
  wire [3:0] _T_333; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296634.4]
  wire  _T_334; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296637.4]
  wire  _T_335; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296638.4]
  wire  _T_336; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296639.4]
  wire  _T_338; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296641.4]
  wire  _T_339; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296642.4]
  wire  _T_340; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296647.4]
  wire  _T_341; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296648.4]
  wire  _T_342; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296649.4]
  wire  _T_344; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296651.4]
  wire  _T_345; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296652.4]
  wire  _T_346; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296657.4]
  reg [3:0] _T_348; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296658.4]
  reg [31:0] _RAND_6;
  wire  _T_350; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296661.4]
  wire  _T_352; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296663.4]
  wire  _T_353; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296664.4]
  wire  _T_354; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296665.4]
  wire  _T_356; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296667.4]
  wire  _T_357; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296668.4]
  wire [3:0] _GEN_106; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296669.4]
  wire [3:0] _T_359; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296670.4]
  wire [3:0] _GEN_107; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296671.4]
  wire [4:0] _T_360; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296671.4]
  wire [4:0] _T_361; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296672.4]
  wire [3:0] _T_362; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296673.4]
  wire  _T_363; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296676.4]
  wire  _T_364; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296677.4]
  wire  _T_365; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296678.4]
  wire  _T_367; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296680.4]
  wire  _T_368; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296681.4]
  wire  _T_369; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296686.4]
  wire  _T_370; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296687.4]
  wire  _T_371; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296688.4]
  wire  _T_373; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296690.4]
  wire  _T_374; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296691.4]
  wire  _T_375; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296696.4]
  reg [3:0] _T_377; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296697.4]
  reg [31:0] _RAND_7;
  wire  _T_379; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296700.4]
  wire  _T_381; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296702.4]
  wire  _T_382; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296703.4]
  wire  _T_383; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296704.4]
  wire  _T_385; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296706.4]
  wire  _T_386; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296707.4]
  wire [3:0] _GEN_108; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296708.4]
  wire [3:0] _T_388; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296709.4]
  wire [3:0] _GEN_109; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296710.4]
  wire [4:0] _T_389; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296710.4]
  wire [4:0] _T_390; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296711.4]
  wire [3:0] _T_391; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296712.4]
  wire  _T_392; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296715.4]
  wire  _T_393; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296716.4]
  wire  _T_394; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296717.4]
  wire  _T_396; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296719.4]
  wire  _T_397; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296720.4]
  wire  _T_398; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296725.4]
  wire  _T_399; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296726.4]
  wire  _T_400; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296727.4]
  wire  _T_402; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296729.4]
  wire  _T_403; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296730.4]
  wire  _T_404; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296735.4]
  reg [3:0] _T_406; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296736.4]
  reg [31:0] _RAND_8;
  wire  _T_408; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296739.4]
  wire  _T_410; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296741.4]
  wire  _T_411; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296742.4]
  wire  _T_412; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296743.4]
  wire  _T_414; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296745.4]
  wire  _T_415; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296746.4]
  wire [3:0] _GEN_110; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296747.4]
  wire [3:0] _T_417; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296748.4]
  wire [3:0] _GEN_111; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296749.4]
  wire [4:0] _T_418; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296749.4]
  wire [4:0] _T_419; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296750.4]
  wire [3:0] _T_420; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296751.4]
  wire  _T_421; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296754.4]
  wire  _T_422; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296755.4]
  wire  _T_423; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296756.4]
  wire  _T_425; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296758.4]
  wire  _T_426; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296759.4]
  wire  _T_427; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296764.4]
  wire  _T_428; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296765.4]
  wire  _T_429; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296766.4]
  wire  _T_431; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296768.4]
  wire  _T_432; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296769.4]
  wire  _T_433; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296774.4]
  reg [3:0] _T_435; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296775.4]
  reg [31:0] _RAND_9;
  wire  _T_437; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296778.4]
  wire  _T_439; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296780.4]
  wire  _T_440; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296781.4]
  wire  _T_441; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296782.4]
  wire  _T_443; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296784.4]
  wire  _T_444; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296785.4]
  wire [3:0] _GEN_112; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296786.4]
  wire [3:0] _T_446; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296787.4]
  wire [3:0] _GEN_113; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296788.4]
  wire [4:0] _T_447; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296788.4]
  wire [4:0] _T_448; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296789.4]
  wire [3:0] _T_449; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296790.4]
  wire  _T_450; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296793.4]
  wire  _T_451; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296794.4]
  wire  _T_452; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296795.4]
  wire  _T_454; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296797.4]
  wire  _T_455; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296798.4]
  wire  _T_456; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296803.4]
  wire  _T_457; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296804.4]
  wire  _T_458; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296805.4]
  wire  _T_460; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296807.4]
  wire  _T_461; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296808.4]
  wire  _T_462; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296813.4]
  reg [3:0] _T_464; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296814.4]
  reg [31:0] _RAND_10;
  wire  _T_466; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296817.4]
  wire  _T_468; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296819.4]
  wire  _T_469; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296820.4]
  wire  _T_470; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296821.4]
  wire  _T_472; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296823.4]
  wire  _T_473; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296824.4]
  wire [3:0] _GEN_114; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296825.4]
  wire [3:0] _T_475; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296826.4]
  wire [3:0] _GEN_115; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296827.4]
  wire [4:0] _T_476; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296827.4]
  wire [4:0] _T_477; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296828.4]
  wire [3:0] _T_478; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296829.4]
  wire  _T_479; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296832.4]
  wire  _T_480; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296833.4]
  wire  _T_481; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296834.4]
  wire  _T_483; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296836.4]
  wire  _T_484; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296837.4]
  wire  _T_485; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296842.4]
  wire  _T_486; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296843.4]
  wire  _T_487; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296844.4]
  wire  _T_489; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296846.4]
  wire  _T_490; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296847.4]
  wire  _T_491; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296852.4]
  reg [3:0] _T_493; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296853.4]
  reg [31:0] _RAND_11;
  wire  _T_495; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296856.4]
  wire  _T_497; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296858.4]
  wire  _T_498; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296859.4]
  wire  _T_499; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296860.4]
  wire  _T_501; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296862.4]
  wire  _T_502; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296863.4]
  wire [3:0] _GEN_116; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296864.4]
  wire [3:0] _T_504; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296865.4]
  wire [3:0] _GEN_117; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296866.4]
  wire [4:0] _T_505; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296866.4]
  wire [4:0] _T_506; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296867.4]
  wire [3:0] _T_507; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296868.4]
  wire  _T_508; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296871.4]
  wire  _T_509; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296872.4]
  wire  _T_510; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296873.4]
  wire  _T_512; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296875.4]
  wire  _T_513; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296876.4]
  wire  _T_514; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296881.4]
  wire  _T_515; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296882.4]
  wire  _T_516; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296883.4]
  wire  _T_518; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296885.4]
  wire  _T_519; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296886.4]
  wire  _T_520; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296891.4]
  reg [3:0] _T_522; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296892.4]
  reg [31:0] _RAND_12;
  wire  _T_524; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296895.4]
  wire  _T_526; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296897.4]
  wire  _T_527; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296898.4]
  wire  _T_528; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296899.4]
  wire  _T_530; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296901.4]
  wire  _T_531; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296902.4]
  wire [3:0] _GEN_118; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296903.4]
  wire [3:0] _T_533; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296904.4]
  wire [3:0] _GEN_119; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296905.4]
  wire [4:0] _T_534; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296905.4]
  wire [4:0] _T_535; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296906.4]
  wire [3:0] _T_536; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296907.4]
  wire  _T_537; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296910.4]
  wire  _T_538; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296911.4]
  wire  _T_539; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296912.4]
  wire  _T_541; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296914.4]
  wire  _T_542; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296915.4]
  wire  _T_543; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296920.4]
  wire  _T_544; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296921.4]
  wire  _T_545; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296922.4]
  wire  _T_547; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296924.4]
  wire  _T_548; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296925.4]
  wire  _T_549; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296930.4]
  reg [3:0] _T_551; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296931.4]
  reg [31:0] _RAND_13;
  wire  _T_553; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296934.4]
  wire  _T_555; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296936.4]
  wire  _T_556; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296937.4]
  wire  _T_557; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296938.4]
  wire  _T_559; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296940.4]
  wire  _T_560; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296941.4]
  wire [3:0] _GEN_120; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296942.4]
  wire [3:0] _T_562; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296943.4]
  wire [3:0] _GEN_121; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296944.4]
  wire [4:0] _T_563; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296944.4]
  wire [4:0] _T_564; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296945.4]
  wire [3:0] _T_565; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296946.4]
  wire  _T_566; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296949.4]
  wire  _T_567; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296950.4]
  wire  _T_568; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296951.4]
  wire  _T_570; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296953.4]
  wire  _T_571; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296954.4]
  wire  _T_572; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296959.4]
  wire  _T_573; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296960.4]
  wire  _T_574; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296961.4]
  wire  _T_576; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296963.4]
  wire  _T_577; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296964.4]
  wire  _T_578; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296969.4]
  reg [3:0] _T_580; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296970.4]
  reg [31:0] _RAND_14;
  wire  _T_582; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296973.4]
  wire  _T_584; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296975.4]
  wire  _T_585; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296976.4]
  wire  _T_586; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296977.4]
  wire  _T_588; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296979.4]
  wire  _T_589; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296980.4]
  wire [3:0] _GEN_122; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296981.4]
  wire [3:0] _T_591; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296982.4]
  wire [3:0] _GEN_123; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296983.4]
  wire [4:0] _T_592; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296983.4]
  wire [4:0] _T_593; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296984.4]
  wire [3:0] _T_594; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296985.4]
  wire  _T_595; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296988.4]
  wire  _T_596; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296989.4]
  wire  _T_597; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296990.4]
  wire  _T_599; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296992.4]
  wire  _T_600; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296993.4]
  wire  _T_601; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296998.4]
  wire  _T_602; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296999.4]
  wire  _T_603; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297000.4]
  wire  _T_605; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297002.4]
  wire  _T_606; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297003.4]
  wire  _T_607; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297008.4]
  reg [3:0] _T_609; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297009.4]
  reg [31:0] _RAND_15;
  wire  _T_611; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297012.4]
  wire  _T_613; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297014.4]
  wire  _T_614; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297015.4]
  wire  _T_615; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297016.4]
  wire  _T_617; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297018.4]
  wire  _T_618; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297019.4]
  wire [3:0] _GEN_124; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297020.4]
  wire [3:0] _T_620; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297021.4]
  wire [3:0] _GEN_125; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297022.4]
  wire [4:0] _T_621; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297022.4]
  wire [4:0] _T_622; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297023.4]
  wire [3:0] _T_623; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297024.4]
  wire  _T_624; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297027.4]
  wire  _T_625; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297028.4]
  wire  _T_626; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297029.4]
  wire  _T_628; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297031.4]
  wire  _T_629; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297032.4]
  wire  _T_630; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297037.4]
  wire  _T_631; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297038.4]
  wire  _T_632; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297039.4]
  wire  _T_634; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297041.4]
  wire  _T_635; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297042.4]
  wire  _T_636; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297047.4]
  reg [3:0] _T_638; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297048.4]
  reg [31:0] _RAND_16;
  wire  _T_640; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297051.4]
  wire  _T_642; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297053.4]
  wire  _T_643; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297054.4]
  wire  _T_644; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297055.4]
  wire  _T_646; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297057.4]
  wire  _T_647; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297058.4]
  wire [3:0] _GEN_126; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297059.4]
  wire [3:0] _T_649; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297060.4]
  wire [3:0] _GEN_127; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297061.4]
  wire [4:0] _T_650; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297061.4]
  wire [4:0] _T_651; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297062.4]
  wire [3:0] _T_652; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297063.4]
  wire  _T_653; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297066.4]
  wire  _T_654; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297067.4]
  wire  _T_655; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297068.4]
  wire  _T_657; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297070.4]
  wire  _T_658; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297071.4]
  wire  _T_659; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297076.4]
  wire  _T_660; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297077.4]
  wire  _T_661; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297078.4]
  wire  _T_663; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297080.4]
  wire  _T_664; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297081.4]
  wire  _T_665; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297086.4]
  reg [3:0] _T_667; // @[Deinterleaver.scala 62:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297087.4]
  reg [31:0] _RAND_17;
  wire  _T_669; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297090.4]
  wire  _T_671; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297092.4]
  wire  _T_672; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297093.4]
  wire  _T_673; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297094.4]
  wire  _T_675; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297096.4]
  wire  _T_676; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297097.4]
  wire [3:0] _GEN_128; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297098.4]
  wire [3:0] _T_678; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297099.4]
  wire [3:0] _GEN_129; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297100.4]
  wire [4:0] _T_679; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297100.4]
  wire [4:0] _T_680; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297101.4]
  wire [3:0] _T_681; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297102.4]
  wire  _T_682; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297105.4]
  wire  _T_683; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297106.4]
  wire  _T_684; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297107.4]
  wire  _T_686; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297109.4]
  wire  _T_687; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297110.4]
  wire  _T_688; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297115.4]
  wire  _T_689; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297116.4]
  wire  _T_690; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297117.4]
  wire  _T_692; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297119.4]
  wire  _T_693; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297120.4]
  wire  _T_694; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297125.4]
  wire [1:0] _T_695; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297126.4]
  wire [1:0] _T_696; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297127.4]
  wire [3:0] _T_697; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297128.4]
  wire [1:0] _T_698; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297129.4]
  wire [1:0] _T_699; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297130.4]
  wire [3:0] _T_700; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297131.4]
  wire [7:0] _T_701; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297132.4]
  wire [1:0] _T_702; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297133.4]
  wire [1:0] _T_703; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297134.4]
  wire [3:0] _T_704; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297135.4]
  wire [1:0] _T_705; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297136.4]
  wire [1:0] _T_706; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297137.4]
  wire [3:0] _T_707; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297138.4]
  wire [7:0] _T_708; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297139.4]
  wire [15:0] _T_709; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297140.4]
  wire [16:0] _GEN_130; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297141.4]
  wire [16:0] _T_710; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297141.4]
  wire [15:0] _T_711; // @[package.scala 194:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297142.4]
  wire [15:0] _T_712; // @[package.scala 194:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297143.4]
  wire [17:0] _GEN_131; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297144.4]
  wire [17:0] _T_713; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297144.4]
  wire [15:0] _T_714; // @[package.scala 194:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297145.4]
  wire [15:0] _T_715; // @[package.scala 194:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297146.4]
  wire [19:0] _GEN_132; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297147.4]
  wire [19:0] _T_716; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297147.4]
  wire [15:0] _T_717; // @[package.scala 194:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297148.4]
  wire [15:0] _T_718; // @[package.scala 194:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297149.4]
  wire [23:0] _GEN_133; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297150.4]
  wire [23:0] _T_719; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297150.4]
  wire [15:0] _T_720; // @[package.scala 194:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297151.4]
  wire [15:0] _T_721; // @[package.scala 194:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297152.4]
  wire [16:0] _GEN_134; // @[Deinterleaver.scala 76:51:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297154.4]
  wire [16:0] _T_723; // @[Deinterleaver.scala 76:51:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297154.4]
  wire [16:0] _T_724; // @[Deinterleaver.scala 76:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297155.4]
  wire [16:0] _T_725; // @[Deinterleaver.scala 76:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297156.4]
  wire  _T_726; // @[Deinterleaver.scala 77:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297157.4]
  wire  _T_728; // @[Deinterleaver.scala 77:39:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297159.4]
  wire  _T_729; // @[Deinterleaver.scala 77:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297160.4]
  wire  _T_730; // @[Deinterleaver.scala 78:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297162.6]
  wire  _T_731; // @[OneHot.scala 26:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297164.6]
  wire [15:0] _T_732; // @[OneHot.scala 27:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297165.6]
  wire [15:0] _GEN_136; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297167.6]
  wire [15:0] _T_734; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297167.6]
  wire [7:0] _T_735; // @[OneHot.scala 26:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297168.6]
  wire [7:0] _T_736; // @[OneHot.scala 27:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297169.6]
  wire  _T_737; // @[OneHot.scala 28:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297170.6]
  wire [7:0] _T_738; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297171.6]
  wire [3:0] _T_739; // @[OneHot.scala 26:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297172.6]
  wire [3:0] _T_740; // @[OneHot.scala 27:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297173.6]
  wire  _T_741; // @[OneHot.scala 28:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297174.6]
  wire [3:0] _T_742; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297175.6]
  wire [1:0] _T_743; // @[OneHot.scala 26:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297176.6]
  wire [1:0] _T_744; // @[OneHot.scala 27:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297177.6]
  wire  _T_745; // @[OneHot.scala 28:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297178.6]
  wire [1:0] _T_746; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297179.6]
  wire  _T_747; // @[CircuitMath.scala 30:8:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297180.6]
  wire [1:0] _T_748; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297181.6]
  wire [2:0] _T_749; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297182.6]
  wire [3:0] _T_750; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297183.6]
  wire [4:0] _T_751; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297184.6]
  wire [4:0] _GEN_1; // @[Deinterleaver.scala 77:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297161.4]
  wire [3:0] _T_755_0_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  wire [63:0] _T_755_0_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  wire [1:0] _T_755_0_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  wire [12:0] _T_755_0_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  wire [3:0] _T_755_1_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  wire [3:0] _GEN_7; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_1_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  wire [63:0] _GEN_8; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_1_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  wire [1:0] _GEN_9; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_1_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  wire [12:0] _GEN_10; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_2_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  wire [3:0] _GEN_12; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_2_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  wire [63:0] _GEN_13; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_2_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  wire [1:0] _GEN_14; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_2_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  wire [12:0] _GEN_15; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_3_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  wire [3:0] _GEN_17; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_3_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  wire [63:0] _GEN_18; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_3_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  wire [1:0] _GEN_19; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_3_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  wire [12:0] _GEN_20; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_4_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  wire [3:0] _GEN_22; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_4_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  wire [63:0] _GEN_23; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_4_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  wire [1:0] _GEN_24; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_4_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  wire [12:0] _GEN_25; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_5_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  wire [3:0] _GEN_27; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_5_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  wire [63:0] _GEN_28; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_5_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  wire [1:0] _GEN_29; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_5_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  wire [12:0] _GEN_30; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_6_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  wire [3:0] _GEN_32; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_6_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  wire [63:0] _GEN_33; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_6_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  wire [1:0] _GEN_34; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_6_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  wire [12:0] _GEN_35; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_7_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  wire [3:0] _GEN_37; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_7_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  wire [63:0] _GEN_38; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_7_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  wire [1:0] _GEN_39; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_7_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  wire [12:0] _GEN_40; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_8_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  wire [3:0] _GEN_42; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_8_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  wire [63:0] _GEN_43; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_8_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  wire [1:0] _GEN_44; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_8_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  wire [12:0] _GEN_45; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_9_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  wire [3:0] _GEN_47; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_9_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  wire [63:0] _GEN_48; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_9_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  wire [1:0] _GEN_49; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_9_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  wire [12:0] _GEN_50; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_10_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  wire [3:0] _GEN_52; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_10_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  wire [63:0] _GEN_53; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_10_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  wire [1:0] _GEN_54; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_10_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  wire [12:0] _GEN_55; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_11_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  wire [3:0] _GEN_57; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_11_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  wire [63:0] _GEN_58; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_11_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  wire [1:0] _GEN_59; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_11_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  wire [12:0] _GEN_60; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_12_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  wire [3:0] _GEN_62; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_12_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  wire [63:0] _GEN_63; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_12_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  wire [1:0] _GEN_64; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_12_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  wire [12:0] _GEN_65; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_13_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  wire [3:0] _GEN_67; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_13_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  wire [63:0] _GEN_68; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_13_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  wire [1:0] _GEN_69; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_13_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  wire [12:0] _GEN_70; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_14_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  wire [3:0] _GEN_72; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [63:0] _T_755_14_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  wire [63:0] _GEN_73; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [1:0] _T_755_14_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  wire [1:0] _GEN_74; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [12:0] _T_755_14_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  wire [12:0] _GEN_75; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  wire [3:0] _T_755_15_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  wire [63:0] _T_755_15_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  wire [1:0] _T_755_15_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  wire [12:0] _T_755_15_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  Queue_46 Queue ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296430.4]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_resp(Queue_io_enq_bits_resp),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_resp(Queue_io_deq_bits_resp),
    .io_deq_bits_user(Queue_io_deq_bits_user),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_46 Queue_1 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296434.4]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_resp(Queue_1_io_enq_bits_resp),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_resp(Queue_1_io_deq_bits_resp),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_46 Queue_2 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296438.4]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_enq_bits_user(Queue_2_io_enq_bits_user),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp),
    .io_deq_bits_user(Queue_2_io_deq_bits_user),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  Queue_46 Queue_3 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296442.4]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_data(Queue_3_io_enq_bits_data),
    .io_enq_bits_resp(Queue_3_io_enq_bits_resp),
    .io_enq_bits_user(Queue_3_io_enq_bits_user),
    .io_enq_bits_last(Queue_3_io_enq_bits_last),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_data(Queue_3_io_deq_bits_data),
    .io_deq_bits_resp(Queue_3_io_deq_bits_resp),
    .io_deq_bits_user(Queue_3_io_deq_bits_user),
    .io_deq_bits_last(Queue_3_io_deq_bits_last)
  );
  Queue_46 Queue_4 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296446.4]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_user(Queue_4_io_enq_bits_user),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_user(Queue_4_io_deq_bits_user),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  Queue_46 Queue_5 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296450.4]
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits_id(Queue_5_io_enq_bits_id),
    .io_enq_bits_data(Queue_5_io_enq_bits_data),
    .io_enq_bits_resp(Queue_5_io_enq_bits_resp),
    .io_enq_bits_user(Queue_5_io_enq_bits_user),
    .io_enq_bits_last(Queue_5_io_enq_bits_last),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits_id(Queue_5_io_deq_bits_id),
    .io_deq_bits_data(Queue_5_io_deq_bits_data),
    .io_deq_bits_resp(Queue_5_io_deq_bits_resp),
    .io_deq_bits_user(Queue_5_io_deq_bits_user),
    .io_deq_bits_last(Queue_5_io_deq_bits_last)
  );
  Queue_46 Queue_6 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296454.4]
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits_id(Queue_6_io_enq_bits_id),
    .io_enq_bits_data(Queue_6_io_enq_bits_data),
    .io_enq_bits_resp(Queue_6_io_enq_bits_resp),
    .io_enq_bits_user(Queue_6_io_enq_bits_user),
    .io_enq_bits_last(Queue_6_io_enq_bits_last),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits_id(Queue_6_io_deq_bits_id),
    .io_deq_bits_data(Queue_6_io_deq_bits_data),
    .io_deq_bits_resp(Queue_6_io_deq_bits_resp),
    .io_deq_bits_user(Queue_6_io_deq_bits_user),
    .io_deq_bits_last(Queue_6_io_deq_bits_last)
  );
  Queue_46 Queue_7 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296458.4]
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits_id(Queue_7_io_enq_bits_id),
    .io_enq_bits_data(Queue_7_io_enq_bits_data),
    .io_enq_bits_resp(Queue_7_io_enq_bits_resp),
    .io_enq_bits_user(Queue_7_io_enq_bits_user),
    .io_enq_bits_last(Queue_7_io_enq_bits_last),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits_id(Queue_7_io_deq_bits_id),
    .io_deq_bits_data(Queue_7_io_deq_bits_data),
    .io_deq_bits_resp(Queue_7_io_deq_bits_resp),
    .io_deq_bits_user(Queue_7_io_deq_bits_user),
    .io_deq_bits_last(Queue_7_io_deq_bits_last)
  );
  Queue_46 Queue_8 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296462.4]
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits_id(Queue_8_io_enq_bits_id),
    .io_enq_bits_data(Queue_8_io_enq_bits_data),
    .io_enq_bits_resp(Queue_8_io_enq_bits_resp),
    .io_enq_bits_user(Queue_8_io_enq_bits_user),
    .io_enq_bits_last(Queue_8_io_enq_bits_last),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits_id(Queue_8_io_deq_bits_id),
    .io_deq_bits_data(Queue_8_io_deq_bits_data),
    .io_deq_bits_resp(Queue_8_io_deq_bits_resp),
    .io_deq_bits_user(Queue_8_io_deq_bits_user),
    .io_deq_bits_last(Queue_8_io_deq_bits_last)
  );
  Queue_46 Queue_9 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296466.4]
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits_id(Queue_9_io_enq_bits_id),
    .io_enq_bits_data(Queue_9_io_enq_bits_data),
    .io_enq_bits_resp(Queue_9_io_enq_bits_resp),
    .io_enq_bits_user(Queue_9_io_enq_bits_user),
    .io_enq_bits_last(Queue_9_io_enq_bits_last),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits_id(Queue_9_io_deq_bits_id),
    .io_deq_bits_data(Queue_9_io_deq_bits_data),
    .io_deq_bits_resp(Queue_9_io_deq_bits_resp),
    .io_deq_bits_user(Queue_9_io_deq_bits_user),
    .io_deq_bits_last(Queue_9_io_deq_bits_last)
  );
  Queue_46 Queue_10 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296470.4]
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits_id(Queue_10_io_enq_bits_id),
    .io_enq_bits_data(Queue_10_io_enq_bits_data),
    .io_enq_bits_resp(Queue_10_io_enq_bits_resp),
    .io_enq_bits_user(Queue_10_io_enq_bits_user),
    .io_enq_bits_last(Queue_10_io_enq_bits_last),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits_id(Queue_10_io_deq_bits_id),
    .io_deq_bits_data(Queue_10_io_deq_bits_data),
    .io_deq_bits_resp(Queue_10_io_deq_bits_resp),
    .io_deq_bits_user(Queue_10_io_deq_bits_user),
    .io_deq_bits_last(Queue_10_io_deq_bits_last)
  );
  Queue_46 Queue_11 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296474.4]
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits_id(Queue_11_io_enq_bits_id),
    .io_enq_bits_data(Queue_11_io_enq_bits_data),
    .io_enq_bits_resp(Queue_11_io_enq_bits_resp),
    .io_enq_bits_user(Queue_11_io_enq_bits_user),
    .io_enq_bits_last(Queue_11_io_enq_bits_last),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits_id(Queue_11_io_deq_bits_id),
    .io_deq_bits_data(Queue_11_io_deq_bits_data),
    .io_deq_bits_resp(Queue_11_io_deq_bits_resp),
    .io_deq_bits_user(Queue_11_io_deq_bits_user),
    .io_deq_bits_last(Queue_11_io_deq_bits_last)
  );
  Queue_46 Queue_12 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296478.4]
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits_id(Queue_12_io_enq_bits_id),
    .io_enq_bits_data(Queue_12_io_enq_bits_data),
    .io_enq_bits_resp(Queue_12_io_enq_bits_resp),
    .io_enq_bits_user(Queue_12_io_enq_bits_user),
    .io_enq_bits_last(Queue_12_io_enq_bits_last),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits_id(Queue_12_io_deq_bits_id),
    .io_deq_bits_data(Queue_12_io_deq_bits_data),
    .io_deq_bits_resp(Queue_12_io_deq_bits_resp),
    .io_deq_bits_user(Queue_12_io_deq_bits_user),
    .io_deq_bits_last(Queue_12_io_deq_bits_last)
  );
  Queue_46 Queue_13 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296482.4]
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits_id(Queue_13_io_enq_bits_id),
    .io_enq_bits_data(Queue_13_io_enq_bits_data),
    .io_enq_bits_resp(Queue_13_io_enq_bits_resp),
    .io_enq_bits_user(Queue_13_io_enq_bits_user),
    .io_enq_bits_last(Queue_13_io_enq_bits_last),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits_id(Queue_13_io_deq_bits_id),
    .io_deq_bits_data(Queue_13_io_deq_bits_data),
    .io_deq_bits_resp(Queue_13_io_deq_bits_resp),
    .io_deq_bits_user(Queue_13_io_deq_bits_user),
    .io_deq_bits_last(Queue_13_io_deq_bits_last)
  );
  Queue_46 Queue_14 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296486.4]
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits_id(Queue_14_io_enq_bits_id),
    .io_enq_bits_data(Queue_14_io_enq_bits_data),
    .io_enq_bits_resp(Queue_14_io_enq_bits_resp),
    .io_enq_bits_user(Queue_14_io_enq_bits_user),
    .io_enq_bits_last(Queue_14_io_enq_bits_last),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits_id(Queue_14_io_deq_bits_id),
    .io_deq_bits_data(Queue_14_io_deq_bits_data),
    .io_deq_bits_resp(Queue_14_io_deq_bits_resp),
    .io_deq_bits_user(Queue_14_io_deq_bits_user),
    .io_deq_bits_last(Queue_14_io_deq_bits_last)
  );
  Queue_46 Queue_15 ( // @[Deinterleaver.scala 43:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296490.4]
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits_id(Queue_15_io_enq_bits_id),
    .io_enq_bits_data(Queue_15_io_enq_bits_data),
    .io_enq_bits_resp(Queue_15_io_enq_bits_resp),
    .io_enq_bits_user(Queue_15_io_enq_bits_user),
    .io_enq_bits_last(Queue_15_io_enq_bits_last),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits_id(Queue_15_io_deq_bits_id),
    .io_deq_bits_data(Queue_15_io_deq_bits_data),
    .io_deq_bits_resp(Queue_15_io_deq_bits_resp),
    .io_deq_bits_user(Queue_15_io_deq_bits_user),
    .io_deq_bits_last(Queue_15_io_deq_bits_last)
  );
  assign _T_226 = 16'h1 << _T_224; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296497.4]
  assign _T_229 = 16'h1 << auto_out_r_bits_id; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296500.4]
  assign _T_234 = _T_229[0]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296505.4]
  assign _T_826_15 = Queue_15_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297288.4]
  assign _T_826_14 = Queue_14_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297287.4]
  assign _T_826_13 = Queue_13_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297286.4]
  assign _T_826_12 = Queue_12_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297285.4]
  assign _T_826_11 = Queue_11_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297284.4]
  assign _T_826_10 = Queue_10_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297283.4]
  assign _T_826_9 = Queue_9_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297282.4]
  assign _T_826_8 = Queue_8_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297281.4]
  assign _T_826_7 = Queue_7_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297280.4]
  assign _T_826_6 = Queue_6_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297279.4]
  assign _T_826_5 = Queue_5_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297278.4]
  assign _T_826_4 = Queue_4_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297277.4]
  assign _T_826_3 = Queue_3_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297276.4]
  assign _T_826_2 = Queue_2_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297275.4]
  assign _T_826_1 = Queue_1_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297274.4]
  assign _T_826_0 = Queue_io_enq_ready; // @[Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297271.4 Deinterleaver.scala 90:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297273.4]
  assign _GEN_83 = 4'h1 == auto_out_r_bits_id ? _T_826_1 : _T_826_0; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_84 = 4'h2 == auto_out_r_bits_id ? _T_826_2 : _GEN_83; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_85 = 4'h3 == auto_out_r_bits_id ? _T_826_3 : _GEN_84; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_86 = 4'h4 == auto_out_r_bits_id ? _T_826_4 : _GEN_85; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_87 = 4'h5 == auto_out_r_bits_id ? _T_826_5 : _GEN_86; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_88 = 4'h6 == auto_out_r_bits_id ? _T_826_6 : _GEN_87; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_89 = 4'h7 == auto_out_r_bits_id ? _T_826_7 : _GEN_88; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_90 = 4'h8 == auto_out_r_bits_id ? _T_826_8 : _GEN_89; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_91 = 4'h9 == auto_out_r_bits_id ? _T_826_9 : _GEN_90; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_92 = 4'ha == auto_out_r_bits_id ? _T_826_10 : _GEN_91; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_93 = 4'hb == auto_out_r_bits_id ? _T_826_11 : _GEN_92; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_94 = 4'hc == auto_out_r_bits_id ? _T_826_12 : _GEN_93; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_95 = 4'hd == auto_out_r_bits_id ? _T_826_13 : _GEN_94; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_96 = 4'he == auto_out_r_bits_id ? _T_826_14 : _GEN_95; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _GEN_97 = 4'hf == auto_out_r_bits_id ? _T_826_15 : _GEN_96; // @[Deinterleaver.scala 90:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297289.4]
  assign _T_235 = _GEN_97 & auto_out_r_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296506.4]
  assign _T_236 = _T_234 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296507.4]
  assign _T_237 = _T_236 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296508.4]
  assign _T_238 = _T_226[0]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296509.4]
  assign _T_239 = auto_in_r_ready & _T_222; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296510.4]
  assign _T_240 = _T_238 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296511.4]
  assign _T_755_15_last = Queue_15_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  assign _T_755_14_last = Queue_14_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  assign _T_755_13_last = Queue_13_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  assign _T_755_12_last = Queue_12_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  assign _T_755_11_last = Queue_11_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  assign _T_755_10_last = Queue_10_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  assign _T_755_9_last = Queue_9_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  assign _T_755_8_last = Queue_8_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  assign _T_755_7_last = Queue_7_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  assign _T_755_6_last = Queue_6_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  assign _T_755_5_last = Queue_5_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  assign _T_755_4_last = Queue_4_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  assign _T_755_3_last = Queue_3_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  assign _T_755_2_last = Queue_2_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  assign _T_755_1_last = Queue_1_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  assign _T_755_0_last = Queue_io_deq_bits_last; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  assign _GEN_11 = 4'h1 == _T_224 ? _T_755_1_last : _T_755_0_last; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_16 = 4'h2 == _T_224 ? _T_755_2_last : _GEN_11; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_21 = 4'h3 == _T_224 ? _T_755_3_last : _GEN_16; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_26 = 4'h4 == _T_224 ? _T_755_4_last : _GEN_21; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_31 = 4'h5 == _T_224 ? _T_755_5_last : _GEN_26; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_36 = 4'h6 == _T_224 ? _T_755_6_last : _GEN_31; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_41 = 4'h7 == _T_224 ? _T_755_7_last : _GEN_36; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_46 = 4'h8 == _T_224 ? _T_755_8_last : _GEN_41; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_51 = 4'h9 == _T_224 ? _T_755_9_last : _GEN_46; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_56 = 4'ha == _T_224 ? _T_755_10_last : _GEN_51; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_61 = 4'hb == _T_224 ? _T_755_11_last : _GEN_56; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_66 = 4'hc == _T_224 ? _T_755_12_last : _GEN_61; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_71 = 4'hd == _T_224 ? _T_755_13_last : _GEN_66; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_76 = 4'he == _T_224 ? _T_755_14_last : _GEN_71; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _GEN_81 = 4'hf == _T_224 ? _T_755_15_last : _GEN_76; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_241 = _T_240 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296512.4]
  assign _GEN_98 = {{3'd0}, _T_237}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296513.4]
  assign _T_243 = _T_232 + _GEN_98; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296514.4]
  assign _GEN_99 = {{3'd0}, _T_241}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296515.4]
  assign _T_244 = _T_243 - _GEN_99; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296515.4]
  assign _T_245 = $unsigned(_T_244); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296516.4]
  assign _T_246 = _T_245[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296517.4]
  assign _T_247 = _T_241 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296520.4]
  assign _T_248 = _T_232 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296521.4]
  assign _T_249 = _T_247 | _T_248; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296522.4]
  assign _T_251 = _T_249 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296524.4]
  assign _T_252 = _T_251 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296525.4]
  assign _T_253 = _T_237 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296530.4]
  assign _T_254 = _T_232 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296531.4]
  assign _T_255 = _T_253 | _T_254; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296532.4]
  assign _T_257 = _T_255 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296534.4]
  assign _T_258 = _T_257 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296535.4]
  assign _T_259 = _T_246 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296540.4]
  assign _T_263 = _T_229[1]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296544.4]
  assign _T_265 = _T_263 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296546.4]
  assign _T_266 = _T_265 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296547.4]
  assign _T_267 = _T_226[1]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296548.4]
  assign _T_269 = _T_267 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296550.4]
  assign _T_270 = _T_269 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296551.4]
  assign _GEN_100 = {{3'd0}, _T_266}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296552.4]
  assign _T_272 = _T_261 + _GEN_100; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296553.4]
  assign _GEN_101 = {{3'd0}, _T_270}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296554.4]
  assign _T_273 = _T_272 - _GEN_101; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296554.4]
  assign _T_274 = $unsigned(_T_273); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296555.4]
  assign _T_275 = _T_274[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296556.4]
  assign _T_276 = _T_270 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296559.4]
  assign _T_277 = _T_261 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296560.4]
  assign _T_278 = _T_276 | _T_277; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296561.4]
  assign _T_280 = _T_278 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296563.4]
  assign _T_281 = _T_280 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296564.4]
  assign _T_282 = _T_266 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296569.4]
  assign _T_283 = _T_261 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296570.4]
  assign _T_284 = _T_282 | _T_283; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296571.4]
  assign _T_286 = _T_284 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296573.4]
  assign _T_287 = _T_286 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296574.4]
  assign _T_288 = _T_275 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296579.4]
  assign _T_292 = _T_229[2]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296583.4]
  assign _T_294 = _T_292 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296585.4]
  assign _T_295 = _T_294 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296586.4]
  assign _T_296 = _T_226[2]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296587.4]
  assign _T_298 = _T_296 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296589.4]
  assign _T_299 = _T_298 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296590.4]
  assign _GEN_102 = {{3'd0}, _T_295}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296591.4]
  assign _T_301 = _T_290 + _GEN_102; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296592.4]
  assign _GEN_103 = {{3'd0}, _T_299}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296593.4]
  assign _T_302 = _T_301 - _GEN_103; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296593.4]
  assign _T_303 = $unsigned(_T_302); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296594.4]
  assign _T_304 = _T_303[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296595.4]
  assign _T_305 = _T_299 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296598.4]
  assign _T_306 = _T_290 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296599.4]
  assign _T_307 = _T_305 | _T_306; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296600.4]
  assign _T_309 = _T_307 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296602.4]
  assign _T_310 = _T_309 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296603.4]
  assign _T_311 = _T_295 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296608.4]
  assign _T_312 = _T_290 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296609.4]
  assign _T_313 = _T_311 | _T_312; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296610.4]
  assign _T_315 = _T_313 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296612.4]
  assign _T_316 = _T_315 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296613.4]
  assign _T_317 = _T_304 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296618.4]
  assign _T_321 = _T_229[3]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296622.4]
  assign _T_323 = _T_321 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296624.4]
  assign _T_324 = _T_323 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296625.4]
  assign _T_325 = _T_226[3]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296626.4]
  assign _T_327 = _T_325 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296628.4]
  assign _T_328 = _T_327 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296629.4]
  assign _GEN_104 = {{3'd0}, _T_324}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296630.4]
  assign _T_330 = _T_319 + _GEN_104; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296631.4]
  assign _GEN_105 = {{3'd0}, _T_328}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296632.4]
  assign _T_331 = _T_330 - _GEN_105; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296632.4]
  assign _T_332 = $unsigned(_T_331); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296633.4]
  assign _T_333 = _T_332[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296634.4]
  assign _T_334 = _T_328 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296637.4]
  assign _T_335 = _T_319 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296638.4]
  assign _T_336 = _T_334 | _T_335; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296639.4]
  assign _T_338 = _T_336 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296641.4]
  assign _T_339 = _T_338 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296642.4]
  assign _T_340 = _T_324 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296647.4]
  assign _T_341 = _T_319 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296648.4]
  assign _T_342 = _T_340 | _T_341; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296649.4]
  assign _T_344 = _T_342 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296651.4]
  assign _T_345 = _T_344 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296652.4]
  assign _T_346 = _T_333 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296657.4]
  assign _T_350 = _T_229[4]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296661.4]
  assign _T_352 = _T_350 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296663.4]
  assign _T_353 = _T_352 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296664.4]
  assign _T_354 = _T_226[4]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296665.4]
  assign _T_356 = _T_354 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296667.4]
  assign _T_357 = _T_356 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296668.4]
  assign _GEN_106 = {{3'd0}, _T_353}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296669.4]
  assign _T_359 = _T_348 + _GEN_106; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296670.4]
  assign _GEN_107 = {{3'd0}, _T_357}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296671.4]
  assign _T_360 = _T_359 - _GEN_107; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296671.4]
  assign _T_361 = $unsigned(_T_360); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296672.4]
  assign _T_362 = _T_361[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296673.4]
  assign _T_363 = _T_357 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296676.4]
  assign _T_364 = _T_348 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296677.4]
  assign _T_365 = _T_363 | _T_364; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296678.4]
  assign _T_367 = _T_365 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296680.4]
  assign _T_368 = _T_367 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296681.4]
  assign _T_369 = _T_353 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296686.4]
  assign _T_370 = _T_348 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296687.4]
  assign _T_371 = _T_369 | _T_370; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296688.4]
  assign _T_373 = _T_371 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296690.4]
  assign _T_374 = _T_373 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296691.4]
  assign _T_375 = _T_362 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296696.4]
  assign _T_379 = _T_229[5]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296700.4]
  assign _T_381 = _T_379 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296702.4]
  assign _T_382 = _T_381 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296703.4]
  assign _T_383 = _T_226[5]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296704.4]
  assign _T_385 = _T_383 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296706.4]
  assign _T_386 = _T_385 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296707.4]
  assign _GEN_108 = {{3'd0}, _T_382}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296708.4]
  assign _T_388 = _T_377 + _GEN_108; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296709.4]
  assign _GEN_109 = {{3'd0}, _T_386}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296710.4]
  assign _T_389 = _T_388 - _GEN_109; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296710.4]
  assign _T_390 = $unsigned(_T_389); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296711.4]
  assign _T_391 = _T_390[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296712.4]
  assign _T_392 = _T_386 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296715.4]
  assign _T_393 = _T_377 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296716.4]
  assign _T_394 = _T_392 | _T_393; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296717.4]
  assign _T_396 = _T_394 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296719.4]
  assign _T_397 = _T_396 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296720.4]
  assign _T_398 = _T_382 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296725.4]
  assign _T_399 = _T_377 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296726.4]
  assign _T_400 = _T_398 | _T_399; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296727.4]
  assign _T_402 = _T_400 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296729.4]
  assign _T_403 = _T_402 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296730.4]
  assign _T_404 = _T_391 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296735.4]
  assign _T_408 = _T_229[6]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296739.4]
  assign _T_410 = _T_408 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296741.4]
  assign _T_411 = _T_410 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296742.4]
  assign _T_412 = _T_226[6]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296743.4]
  assign _T_414 = _T_412 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296745.4]
  assign _T_415 = _T_414 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296746.4]
  assign _GEN_110 = {{3'd0}, _T_411}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296747.4]
  assign _T_417 = _T_406 + _GEN_110; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296748.4]
  assign _GEN_111 = {{3'd0}, _T_415}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296749.4]
  assign _T_418 = _T_417 - _GEN_111; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296749.4]
  assign _T_419 = $unsigned(_T_418); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296750.4]
  assign _T_420 = _T_419[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296751.4]
  assign _T_421 = _T_415 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296754.4]
  assign _T_422 = _T_406 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296755.4]
  assign _T_423 = _T_421 | _T_422; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296756.4]
  assign _T_425 = _T_423 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296758.4]
  assign _T_426 = _T_425 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296759.4]
  assign _T_427 = _T_411 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296764.4]
  assign _T_428 = _T_406 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296765.4]
  assign _T_429 = _T_427 | _T_428; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296766.4]
  assign _T_431 = _T_429 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296768.4]
  assign _T_432 = _T_431 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296769.4]
  assign _T_433 = _T_420 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296774.4]
  assign _T_437 = _T_229[7]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296778.4]
  assign _T_439 = _T_437 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296780.4]
  assign _T_440 = _T_439 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296781.4]
  assign _T_441 = _T_226[7]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296782.4]
  assign _T_443 = _T_441 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296784.4]
  assign _T_444 = _T_443 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296785.4]
  assign _GEN_112 = {{3'd0}, _T_440}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296786.4]
  assign _T_446 = _T_435 + _GEN_112; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296787.4]
  assign _GEN_113 = {{3'd0}, _T_444}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296788.4]
  assign _T_447 = _T_446 - _GEN_113; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296788.4]
  assign _T_448 = $unsigned(_T_447); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296789.4]
  assign _T_449 = _T_448[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296790.4]
  assign _T_450 = _T_444 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296793.4]
  assign _T_451 = _T_435 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296794.4]
  assign _T_452 = _T_450 | _T_451; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296795.4]
  assign _T_454 = _T_452 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296797.4]
  assign _T_455 = _T_454 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296798.4]
  assign _T_456 = _T_440 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296803.4]
  assign _T_457 = _T_435 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296804.4]
  assign _T_458 = _T_456 | _T_457; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296805.4]
  assign _T_460 = _T_458 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296807.4]
  assign _T_461 = _T_460 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296808.4]
  assign _T_462 = _T_449 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296813.4]
  assign _T_466 = _T_229[8]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296817.4]
  assign _T_468 = _T_466 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296819.4]
  assign _T_469 = _T_468 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296820.4]
  assign _T_470 = _T_226[8]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296821.4]
  assign _T_472 = _T_470 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296823.4]
  assign _T_473 = _T_472 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296824.4]
  assign _GEN_114 = {{3'd0}, _T_469}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296825.4]
  assign _T_475 = _T_464 + _GEN_114; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296826.4]
  assign _GEN_115 = {{3'd0}, _T_473}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296827.4]
  assign _T_476 = _T_475 - _GEN_115; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296827.4]
  assign _T_477 = $unsigned(_T_476); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296828.4]
  assign _T_478 = _T_477[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296829.4]
  assign _T_479 = _T_473 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296832.4]
  assign _T_480 = _T_464 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296833.4]
  assign _T_481 = _T_479 | _T_480; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296834.4]
  assign _T_483 = _T_481 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296836.4]
  assign _T_484 = _T_483 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296837.4]
  assign _T_485 = _T_469 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296842.4]
  assign _T_486 = _T_464 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296843.4]
  assign _T_487 = _T_485 | _T_486; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296844.4]
  assign _T_489 = _T_487 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296846.4]
  assign _T_490 = _T_489 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296847.4]
  assign _T_491 = _T_478 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296852.4]
  assign _T_495 = _T_229[9]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296856.4]
  assign _T_497 = _T_495 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296858.4]
  assign _T_498 = _T_497 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296859.4]
  assign _T_499 = _T_226[9]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296860.4]
  assign _T_501 = _T_499 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296862.4]
  assign _T_502 = _T_501 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296863.4]
  assign _GEN_116 = {{3'd0}, _T_498}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296864.4]
  assign _T_504 = _T_493 + _GEN_116; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296865.4]
  assign _GEN_117 = {{3'd0}, _T_502}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296866.4]
  assign _T_505 = _T_504 - _GEN_117; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296866.4]
  assign _T_506 = $unsigned(_T_505); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296867.4]
  assign _T_507 = _T_506[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296868.4]
  assign _T_508 = _T_502 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296871.4]
  assign _T_509 = _T_493 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296872.4]
  assign _T_510 = _T_508 | _T_509; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296873.4]
  assign _T_512 = _T_510 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296875.4]
  assign _T_513 = _T_512 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296876.4]
  assign _T_514 = _T_498 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296881.4]
  assign _T_515 = _T_493 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296882.4]
  assign _T_516 = _T_514 | _T_515; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296883.4]
  assign _T_518 = _T_516 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296885.4]
  assign _T_519 = _T_518 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296886.4]
  assign _T_520 = _T_507 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296891.4]
  assign _T_524 = _T_229[10]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296895.4]
  assign _T_526 = _T_524 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296897.4]
  assign _T_527 = _T_526 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296898.4]
  assign _T_528 = _T_226[10]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296899.4]
  assign _T_530 = _T_528 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296901.4]
  assign _T_531 = _T_530 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296902.4]
  assign _GEN_118 = {{3'd0}, _T_527}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296903.4]
  assign _T_533 = _T_522 + _GEN_118; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296904.4]
  assign _GEN_119 = {{3'd0}, _T_531}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296905.4]
  assign _T_534 = _T_533 - _GEN_119; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296905.4]
  assign _T_535 = $unsigned(_T_534); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296906.4]
  assign _T_536 = _T_535[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296907.4]
  assign _T_537 = _T_531 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296910.4]
  assign _T_538 = _T_522 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296911.4]
  assign _T_539 = _T_537 | _T_538; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296912.4]
  assign _T_541 = _T_539 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296914.4]
  assign _T_542 = _T_541 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296915.4]
  assign _T_543 = _T_527 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296920.4]
  assign _T_544 = _T_522 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296921.4]
  assign _T_545 = _T_543 | _T_544; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296922.4]
  assign _T_547 = _T_545 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296924.4]
  assign _T_548 = _T_547 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296925.4]
  assign _T_549 = _T_536 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296930.4]
  assign _T_553 = _T_229[11]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296934.4]
  assign _T_555 = _T_553 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296936.4]
  assign _T_556 = _T_555 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296937.4]
  assign _T_557 = _T_226[11]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296938.4]
  assign _T_559 = _T_557 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296940.4]
  assign _T_560 = _T_559 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296941.4]
  assign _GEN_120 = {{3'd0}, _T_556}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296942.4]
  assign _T_562 = _T_551 + _GEN_120; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296943.4]
  assign _GEN_121 = {{3'd0}, _T_560}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296944.4]
  assign _T_563 = _T_562 - _GEN_121; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296944.4]
  assign _T_564 = $unsigned(_T_563); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296945.4]
  assign _T_565 = _T_564[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296946.4]
  assign _T_566 = _T_560 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296949.4]
  assign _T_567 = _T_551 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296950.4]
  assign _T_568 = _T_566 | _T_567; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296951.4]
  assign _T_570 = _T_568 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296953.4]
  assign _T_571 = _T_570 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296954.4]
  assign _T_572 = _T_556 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296959.4]
  assign _T_573 = _T_551 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296960.4]
  assign _T_574 = _T_572 | _T_573; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296961.4]
  assign _T_576 = _T_574 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296963.4]
  assign _T_577 = _T_576 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296964.4]
  assign _T_578 = _T_565 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296969.4]
  assign _T_582 = _T_229[12]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296973.4]
  assign _T_584 = _T_582 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296975.4]
  assign _T_585 = _T_584 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296976.4]
  assign _T_586 = _T_226[12]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296977.4]
  assign _T_588 = _T_586 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296979.4]
  assign _T_589 = _T_588 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296980.4]
  assign _GEN_122 = {{3'd0}, _T_585}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296981.4]
  assign _T_591 = _T_580 + _GEN_122; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296982.4]
  assign _GEN_123 = {{3'd0}, _T_589}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296983.4]
  assign _T_592 = _T_591 - _GEN_123; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296983.4]
  assign _T_593 = $unsigned(_T_592); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296984.4]
  assign _T_594 = _T_593[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296985.4]
  assign _T_595 = _T_589 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296988.4]
  assign _T_596 = _T_580 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296989.4]
  assign _T_597 = _T_595 | _T_596; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296990.4]
  assign _T_599 = _T_597 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296992.4]
  assign _T_600 = _T_599 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296993.4]
  assign _T_601 = _T_585 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296998.4]
  assign _T_602 = _T_580 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296999.4]
  assign _T_603 = _T_601 | _T_602; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297000.4]
  assign _T_605 = _T_603 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297002.4]
  assign _T_606 = _T_605 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297003.4]
  assign _T_607 = _T_594 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297008.4]
  assign _T_611 = _T_229[13]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297012.4]
  assign _T_613 = _T_611 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297014.4]
  assign _T_614 = _T_613 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297015.4]
  assign _T_615 = _T_226[13]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297016.4]
  assign _T_617 = _T_615 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297018.4]
  assign _T_618 = _T_617 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297019.4]
  assign _GEN_124 = {{3'd0}, _T_614}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297020.4]
  assign _T_620 = _T_609 + _GEN_124; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297021.4]
  assign _GEN_125 = {{3'd0}, _T_618}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297022.4]
  assign _T_621 = _T_620 - _GEN_125; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297022.4]
  assign _T_622 = $unsigned(_T_621); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297023.4]
  assign _T_623 = _T_622[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297024.4]
  assign _T_624 = _T_618 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297027.4]
  assign _T_625 = _T_609 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297028.4]
  assign _T_626 = _T_624 | _T_625; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297029.4]
  assign _T_628 = _T_626 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297031.4]
  assign _T_629 = _T_628 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297032.4]
  assign _T_630 = _T_614 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297037.4]
  assign _T_631 = _T_609 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297038.4]
  assign _T_632 = _T_630 | _T_631; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297039.4]
  assign _T_634 = _T_632 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297041.4]
  assign _T_635 = _T_634 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297042.4]
  assign _T_636 = _T_623 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297047.4]
  assign _T_640 = _T_229[14]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297051.4]
  assign _T_642 = _T_640 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297053.4]
  assign _T_643 = _T_642 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297054.4]
  assign _T_644 = _T_226[14]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297055.4]
  assign _T_646 = _T_644 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297057.4]
  assign _T_647 = _T_646 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297058.4]
  assign _GEN_126 = {{3'd0}, _T_643}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297059.4]
  assign _T_649 = _T_638 + _GEN_126; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297060.4]
  assign _GEN_127 = {{3'd0}, _T_647}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297061.4]
  assign _T_650 = _T_649 - _GEN_127; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297061.4]
  assign _T_651 = $unsigned(_T_650); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297062.4]
  assign _T_652 = _T_651[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297063.4]
  assign _T_653 = _T_647 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297066.4]
  assign _T_654 = _T_638 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297067.4]
  assign _T_655 = _T_653 | _T_654; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297068.4]
  assign _T_657 = _T_655 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297070.4]
  assign _T_658 = _T_657 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297071.4]
  assign _T_659 = _T_643 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297076.4]
  assign _T_660 = _T_638 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297077.4]
  assign _T_661 = _T_659 | _T_660; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297078.4]
  assign _T_663 = _T_661 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297080.4]
  assign _T_664 = _T_663 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297081.4]
  assign _T_665 = _T_652 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297086.4]
  assign _T_669 = _T_229[15]; // @[Deinterleaver.scala 64:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297090.4]
  assign _T_671 = _T_669 & _T_235; // @[Deinterleaver.scala 64:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297092.4]
  assign _T_672 = _T_671 & auto_out_r_bits_last; // @[Deinterleaver.scala 64:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297093.4]
  assign _T_673 = _T_226[15]; // @[Deinterleaver.scala 65:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297094.4]
  assign _T_675 = _T_673 & _T_239; // @[Deinterleaver.scala 65:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297096.4]
  assign _T_676 = _T_675 & _GEN_81; // @[Deinterleaver.scala 65:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297097.4]
  assign _GEN_128 = {{3'd0}, _T_672}; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297098.4]
  assign _T_678 = _T_667 + _GEN_128; // @[Deinterleaver.scala 66:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297099.4]
  assign _GEN_129 = {{3'd0}, _T_676}; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297100.4]
  assign _T_679 = _T_678 - _GEN_129; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297100.4]
  assign _T_680 = $unsigned(_T_679); // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297101.4]
  assign _T_681 = _T_680[3:0]; // @[Deinterleaver.scala 66:40:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297102.4]
  assign _T_682 = _T_676 == 1'h0; // @[Deinterleaver.scala 69:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297105.4]
  assign _T_683 = _T_667 != 4'h0; // @[Deinterleaver.scala 69:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297106.4]
  assign _T_684 = _T_682 | _T_683; // @[Deinterleaver.scala 69:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297107.4]
  assign _T_686 = _T_684 | reset; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297109.4]
  assign _T_687 = _T_686 == 1'h0; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297110.4]
  assign _T_688 = _T_672 == 1'h0; // @[Deinterleaver.scala 70:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297115.4]
  assign _T_689 = _T_667 != 4'h8; // @[Deinterleaver.scala 70:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297116.4]
  assign _T_690 = _T_688 | _T_689; // @[Deinterleaver.scala 70:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297117.4]
  assign _T_692 = _T_690 | reset; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297119.4]
  assign _T_693 = _T_692 == 1'h0; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297120.4]
  assign _T_694 = _T_681 != 4'h0; // @[Deinterleaver.scala 71:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297125.4]
  assign _T_695 = {_T_288,_T_259}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297126.4]
  assign _T_696 = {_T_346,_T_317}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297127.4]
  assign _T_697 = {_T_696,_T_695}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297128.4]
  assign _T_698 = {_T_404,_T_375}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297129.4]
  assign _T_699 = {_T_462,_T_433}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297130.4]
  assign _T_700 = {_T_699,_T_698}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297131.4]
  assign _T_701 = {_T_700,_T_697}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297132.4]
  assign _T_702 = {_T_520,_T_491}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297133.4]
  assign _T_703 = {_T_578,_T_549}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297134.4]
  assign _T_704 = {_T_703,_T_702}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297135.4]
  assign _T_705 = {_T_636,_T_607}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297136.4]
  assign _T_706 = {_T_694,_T_665}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297137.4]
  assign _T_707 = {_T_706,_T_705}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297138.4]
  assign _T_708 = {_T_707,_T_704}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297139.4]
  assign _T_709 = {_T_708,_T_701}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297140.4]
  assign _GEN_130 = {{1'd0}, _T_709}; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297141.4]
  assign _T_710 = _GEN_130 << 1; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297141.4]
  assign _T_711 = _T_710[15:0]; // @[package.scala 194:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297142.4]
  assign _T_712 = _T_709 | _T_711; // @[package.scala 194:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297143.4]
  assign _GEN_131 = {{2'd0}, _T_712}; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297144.4]
  assign _T_713 = _GEN_131 << 2; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297144.4]
  assign _T_714 = _T_713[15:0]; // @[package.scala 194:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297145.4]
  assign _T_715 = _T_712 | _T_714; // @[package.scala 194:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297146.4]
  assign _GEN_132 = {{4'd0}, _T_715}; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297147.4]
  assign _T_716 = _GEN_132 << 4; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297147.4]
  assign _T_717 = _T_716[15:0]; // @[package.scala 194:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297148.4]
  assign _T_718 = _T_715 | _T_717; // @[package.scala 194:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297149.4]
  assign _GEN_133 = {{8'd0}, _T_718}; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297150.4]
  assign _T_719 = _GEN_133 << 8; // @[package.scala 194:48:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297150.4]
  assign _T_720 = _T_719[15:0]; // @[package.scala 194:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297151.4]
  assign _T_721 = _T_718 | _T_720; // @[package.scala 194:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297152.4]
  assign _GEN_134 = {{1'd0}, _T_721}; // @[Deinterleaver.scala 76:51:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297154.4]
  assign _T_723 = _GEN_134 << 1; // @[Deinterleaver.scala 76:51:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297154.4]
  assign _T_724 = ~ _T_723; // @[Deinterleaver.scala 76:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297155.4]
  assign _T_725 = _GEN_130 & _T_724; // @[Deinterleaver.scala 76:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297156.4]
  assign _T_726 = _T_222 == 1'h0; // @[Deinterleaver.scala 77:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297157.4]
  assign _T_728 = _T_239 & _GEN_81; // @[Deinterleaver.scala 77:39:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297159.4]
  assign _T_729 = _T_726 | _T_728; // @[Deinterleaver.scala 77:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297160.4]
  assign _T_730 = _T_709 != 16'h0; // @[Deinterleaver.scala 78:29:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297162.6]
  assign _T_731 = _T_725[16]; // @[OneHot.scala 26:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297164.6]
  assign _T_732 = _T_725[15:0]; // @[OneHot.scala 27:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297165.6]
  assign _GEN_136 = {{15'd0}, _T_731}; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297167.6]
  assign _T_734 = _GEN_136 | _T_732; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297167.6]
  assign _T_735 = _T_734[15:8]; // @[OneHot.scala 26:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297168.6]
  assign _T_736 = _T_734[7:0]; // @[OneHot.scala 27:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297169.6]
  assign _T_737 = _T_735 != 8'h0; // @[OneHot.scala 28:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297170.6]
  assign _T_738 = _T_735 | _T_736; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297171.6]
  assign _T_739 = _T_738[7:4]; // @[OneHot.scala 26:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297172.6]
  assign _T_740 = _T_738[3:0]; // @[OneHot.scala 27:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297173.6]
  assign _T_741 = _T_739 != 4'h0; // @[OneHot.scala 28:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297174.6]
  assign _T_742 = _T_739 | _T_740; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297175.6]
  assign _T_743 = _T_742[3:2]; // @[OneHot.scala 26:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297176.6]
  assign _T_744 = _T_742[1:0]; // @[OneHot.scala 27:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297177.6]
  assign _T_745 = _T_743 != 2'h0; // @[OneHot.scala 28:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297178.6]
  assign _T_746 = _T_743 | _T_744; // @[OneHot.scala 28:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297179.6]
  assign _T_747 = _T_746[1]; // @[CircuitMath.scala 30:8:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297180.6]
  assign _T_748 = {_T_745,_T_747}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297181.6]
  assign _T_749 = {_T_741,_T_748}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297182.6]
  assign _T_750 = {_T_737,_T_749}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297183.6]
  assign _T_751 = {_T_731,_T_750}; // @[Cat.scala 30:58:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297184.6]
  assign _GEN_1 = _T_729 ? _T_751 : {{1'd0}, _T_224}; // @[Deinterleaver.scala 77:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297161.4]
  assign _T_755_0_id = Queue_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  assign _T_755_0_data = Queue_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  assign _T_755_0_resp = Queue_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  assign _T_755_0_user = Queue_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297190.4]
  assign _T_755_1_id = Queue_1_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  assign _GEN_7 = 4'h1 == _T_224 ? _T_755_1_id : _T_755_0_id; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_1_data = Queue_1_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  assign _GEN_8 = 4'h1 == _T_224 ? _T_755_1_data : _T_755_0_data; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_1_resp = Queue_1_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  assign _GEN_9 = 4'h1 == _T_224 ? _T_755_1_resp : _T_755_0_resp; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_1_user = Queue_1_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297191.4]
  assign _GEN_10 = 4'h1 == _T_224 ? _T_755_1_user : _T_755_0_user; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_2_id = Queue_2_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  assign _GEN_12 = 4'h2 == _T_224 ? _T_755_2_id : _GEN_7; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_2_data = Queue_2_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  assign _GEN_13 = 4'h2 == _T_224 ? _T_755_2_data : _GEN_8; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_2_resp = Queue_2_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  assign _GEN_14 = 4'h2 == _T_224 ? _T_755_2_resp : _GEN_9; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_2_user = Queue_2_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297192.4]
  assign _GEN_15 = 4'h2 == _T_224 ? _T_755_2_user : _GEN_10; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_3_id = Queue_3_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  assign _GEN_17 = 4'h3 == _T_224 ? _T_755_3_id : _GEN_12; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_3_data = Queue_3_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  assign _GEN_18 = 4'h3 == _T_224 ? _T_755_3_data : _GEN_13; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_3_resp = Queue_3_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  assign _GEN_19 = 4'h3 == _T_224 ? _T_755_3_resp : _GEN_14; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_3_user = Queue_3_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297193.4]
  assign _GEN_20 = 4'h3 == _T_224 ? _T_755_3_user : _GEN_15; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_4_id = Queue_4_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  assign _GEN_22 = 4'h4 == _T_224 ? _T_755_4_id : _GEN_17; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_4_data = Queue_4_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  assign _GEN_23 = 4'h4 == _T_224 ? _T_755_4_data : _GEN_18; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_4_resp = Queue_4_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  assign _GEN_24 = 4'h4 == _T_224 ? _T_755_4_resp : _GEN_19; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_4_user = Queue_4_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297194.4]
  assign _GEN_25 = 4'h4 == _T_224 ? _T_755_4_user : _GEN_20; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_5_id = Queue_5_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  assign _GEN_27 = 4'h5 == _T_224 ? _T_755_5_id : _GEN_22; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_5_data = Queue_5_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  assign _GEN_28 = 4'h5 == _T_224 ? _T_755_5_data : _GEN_23; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_5_resp = Queue_5_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  assign _GEN_29 = 4'h5 == _T_224 ? _T_755_5_resp : _GEN_24; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_5_user = Queue_5_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297195.4]
  assign _GEN_30 = 4'h5 == _T_224 ? _T_755_5_user : _GEN_25; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_6_id = Queue_6_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  assign _GEN_32 = 4'h6 == _T_224 ? _T_755_6_id : _GEN_27; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_6_data = Queue_6_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  assign _GEN_33 = 4'h6 == _T_224 ? _T_755_6_data : _GEN_28; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_6_resp = Queue_6_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  assign _GEN_34 = 4'h6 == _T_224 ? _T_755_6_resp : _GEN_29; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_6_user = Queue_6_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297196.4]
  assign _GEN_35 = 4'h6 == _T_224 ? _T_755_6_user : _GEN_30; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_7_id = Queue_7_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  assign _GEN_37 = 4'h7 == _T_224 ? _T_755_7_id : _GEN_32; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_7_data = Queue_7_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  assign _GEN_38 = 4'h7 == _T_224 ? _T_755_7_data : _GEN_33; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_7_resp = Queue_7_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  assign _GEN_39 = 4'h7 == _T_224 ? _T_755_7_resp : _GEN_34; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_7_user = Queue_7_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297197.4]
  assign _GEN_40 = 4'h7 == _T_224 ? _T_755_7_user : _GEN_35; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_8_id = Queue_8_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  assign _GEN_42 = 4'h8 == _T_224 ? _T_755_8_id : _GEN_37; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_8_data = Queue_8_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  assign _GEN_43 = 4'h8 == _T_224 ? _T_755_8_data : _GEN_38; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_8_resp = Queue_8_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  assign _GEN_44 = 4'h8 == _T_224 ? _T_755_8_resp : _GEN_39; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_8_user = Queue_8_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297198.4]
  assign _GEN_45 = 4'h8 == _T_224 ? _T_755_8_user : _GEN_40; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_9_id = Queue_9_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  assign _GEN_47 = 4'h9 == _T_224 ? _T_755_9_id : _GEN_42; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_9_data = Queue_9_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  assign _GEN_48 = 4'h9 == _T_224 ? _T_755_9_data : _GEN_43; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_9_resp = Queue_9_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  assign _GEN_49 = 4'h9 == _T_224 ? _T_755_9_resp : _GEN_44; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_9_user = Queue_9_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297199.4]
  assign _GEN_50 = 4'h9 == _T_224 ? _T_755_9_user : _GEN_45; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_10_id = Queue_10_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  assign _GEN_52 = 4'ha == _T_224 ? _T_755_10_id : _GEN_47; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_10_data = Queue_10_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  assign _GEN_53 = 4'ha == _T_224 ? _T_755_10_data : _GEN_48; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_10_resp = Queue_10_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  assign _GEN_54 = 4'ha == _T_224 ? _T_755_10_resp : _GEN_49; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_10_user = Queue_10_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297200.4]
  assign _GEN_55 = 4'ha == _T_224 ? _T_755_10_user : _GEN_50; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_11_id = Queue_11_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  assign _GEN_57 = 4'hb == _T_224 ? _T_755_11_id : _GEN_52; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_11_data = Queue_11_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  assign _GEN_58 = 4'hb == _T_224 ? _T_755_11_data : _GEN_53; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_11_resp = Queue_11_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  assign _GEN_59 = 4'hb == _T_224 ? _T_755_11_resp : _GEN_54; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_11_user = Queue_11_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297201.4]
  assign _GEN_60 = 4'hb == _T_224 ? _T_755_11_user : _GEN_55; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_12_id = Queue_12_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  assign _GEN_62 = 4'hc == _T_224 ? _T_755_12_id : _GEN_57; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_12_data = Queue_12_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  assign _GEN_63 = 4'hc == _T_224 ? _T_755_12_data : _GEN_58; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_12_resp = Queue_12_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  assign _GEN_64 = 4'hc == _T_224 ? _T_755_12_resp : _GEN_59; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_12_user = Queue_12_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297202.4]
  assign _GEN_65 = 4'hc == _T_224 ? _T_755_12_user : _GEN_60; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_13_id = Queue_13_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  assign _GEN_67 = 4'hd == _T_224 ? _T_755_13_id : _GEN_62; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_13_data = Queue_13_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  assign _GEN_68 = 4'hd == _T_224 ? _T_755_13_data : _GEN_63; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_13_resp = Queue_13_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  assign _GEN_69 = 4'hd == _T_224 ? _T_755_13_resp : _GEN_64; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_13_user = Queue_13_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297203.4]
  assign _GEN_70 = 4'hd == _T_224 ? _T_755_13_user : _GEN_65; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_14_id = Queue_14_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  assign _GEN_72 = 4'he == _T_224 ? _T_755_14_id : _GEN_67; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_14_data = Queue_14_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  assign _GEN_73 = 4'he == _T_224 ? _T_755_14_data : _GEN_68; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_14_resp = Queue_14_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  assign _GEN_74 = 4'he == _T_224 ? _T_755_14_resp : _GEN_69; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_14_user = Queue_14_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297204.4]
  assign _GEN_75 = 4'he == _T_224 ? _T_755_14_user : _GEN_70; // @[Deinterleaver.scala 84:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297206.4]
  assign _T_755_15_id = Queue_15_io_deq_bits_id; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  assign _T_755_15_data = Queue_15_io_deq_bits_data; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  assign _T_755_15_resp = Queue_15_io_deq_bits_resp; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  assign _T_755_15_user = Queue_15_io_deq_bits_user; // @[Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297188.4 Deinterleaver.scala 84:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297205.4]
  assign auto_in_aw_ready = auto_out_aw_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_b_bits_user = auto_out_b_bits_user; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_r_valid = _T_222; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_r_bits_id = 4'hf == _T_224 ? _T_755_15_id : _GEN_72; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_r_bits_data = 4'hf == _T_224 ? _T_755_15_data : _GEN_73; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_r_bits_resp = 4'hf == _T_224 ? _T_755_15_resp : _GEN_74; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_r_bits_user = 4'hf == _T_224 ? _T_755_15_user : _GEN_75; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_in_r_bits_last = 4'hf == _T_224 ? _T_755_15_last : _GEN_76; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296425.4]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_aw_bits_user = auto_in_aw_bits_user; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_ar_bits_user = auto_in_ar_bits_user; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign auto_out_r_ready = 4'hf == auto_out_r_bits_id ? _T_826_15 : _GEN_96; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296424.4]
  assign Queue_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296432.4]
  assign Queue_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296433.4]
  assign Queue_io_enq_valid = _T_234 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297307.4]
  assign Queue_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297308.4]
  assign Queue_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297308.4]
  assign Queue_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297308.4]
  assign Queue_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297308.4]
  assign Queue_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297308.4]
  assign Queue_io_deq_ready = _T_238 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297225.4]
  assign Queue_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296436.4]
  assign Queue_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296437.4]
  assign Queue_1_io_enq_valid = _T_263 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297310.4]
  assign Queue_1_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297311.4]
  assign Queue_1_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297311.4]
  assign Queue_1_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297311.4]
  assign Queue_1_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297311.4]
  assign Queue_1_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297311.4]
  assign Queue_1_io_deq_ready = _T_267 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297228.4]
  assign Queue_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296440.4]
  assign Queue_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296441.4]
  assign Queue_2_io_enq_valid = _T_292 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297313.4]
  assign Queue_2_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297314.4]
  assign Queue_2_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297314.4]
  assign Queue_2_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297314.4]
  assign Queue_2_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297314.4]
  assign Queue_2_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297314.4]
  assign Queue_2_io_deq_ready = _T_296 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297231.4]
  assign Queue_3_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296444.4]
  assign Queue_3_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296445.4]
  assign Queue_3_io_enq_valid = _T_321 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297316.4]
  assign Queue_3_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297317.4]
  assign Queue_3_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297317.4]
  assign Queue_3_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297317.4]
  assign Queue_3_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297317.4]
  assign Queue_3_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297317.4]
  assign Queue_3_io_deq_ready = _T_325 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297234.4]
  assign Queue_4_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296448.4]
  assign Queue_4_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296449.4]
  assign Queue_4_io_enq_valid = _T_350 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297319.4]
  assign Queue_4_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297320.4]
  assign Queue_4_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297320.4]
  assign Queue_4_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297320.4]
  assign Queue_4_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297320.4]
  assign Queue_4_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297320.4]
  assign Queue_4_io_deq_ready = _T_354 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297237.4]
  assign Queue_5_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296452.4]
  assign Queue_5_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296453.4]
  assign Queue_5_io_enq_valid = _T_379 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297322.4]
  assign Queue_5_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297323.4]
  assign Queue_5_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297323.4]
  assign Queue_5_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297323.4]
  assign Queue_5_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297323.4]
  assign Queue_5_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297323.4]
  assign Queue_5_io_deq_ready = _T_383 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297240.4]
  assign Queue_6_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296456.4]
  assign Queue_6_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296457.4]
  assign Queue_6_io_enq_valid = _T_408 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297325.4]
  assign Queue_6_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297326.4]
  assign Queue_6_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297326.4]
  assign Queue_6_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297326.4]
  assign Queue_6_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297326.4]
  assign Queue_6_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297326.4]
  assign Queue_6_io_deq_ready = _T_412 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297243.4]
  assign Queue_7_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296460.4]
  assign Queue_7_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296461.4]
  assign Queue_7_io_enq_valid = _T_437 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297328.4]
  assign Queue_7_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297329.4]
  assign Queue_7_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297329.4]
  assign Queue_7_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297329.4]
  assign Queue_7_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297329.4]
  assign Queue_7_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297329.4]
  assign Queue_7_io_deq_ready = _T_441 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297246.4]
  assign Queue_8_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296464.4]
  assign Queue_8_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296465.4]
  assign Queue_8_io_enq_valid = _T_466 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297331.4]
  assign Queue_8_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297332.4]
  assign Queue_8_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297332.4]
  assign Queue_8_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297332.4]
  assign Queue_8_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297332.4]
  assign Queue_8_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297332.4]
  assign Queue_8_io_deq_ready = _T_470 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297249.4]
  assign Queue_9_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296468.4]
  assign Queue_9_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296469.4]
  assign Queue_9_io_enq_valid = _T_495 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297334.4]
  assign Queue_9_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297335.4]
  assign Queue_9_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297335.4]
  assign Queue_9_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297335.4]
  assign Queue_9_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297335.4]
  assign Queue_9_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297335.4]
  assign Queue_9_io_deq_ready = _T_499 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297252.4]
  assign Queue_10_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296472.4]
  assign Queue_10_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296473.4]
  assign Queue_10_io_enq_valid = _T_524 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297337.4]
  assign Queue_10_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297338.4]
  assign Queue_10_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297338.4]
  assign Queue_10_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297338.4]
  assign Queue_10_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297338.4]
  assign Queue_10_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297338.4]
  assign Queue_10_io_deq_ready = _T_528 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297255.4]
  assign Queue_11_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296476.4]
  assign Queue_11_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296477.4]
  assign Queue_11_io_enq_valid = _T_553 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297340.4]
  assign Queue_11_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297341.4]
  assign Queue_11_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297341.4]
  assign Queue_11_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297341.4]
  assign Queue_11_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297341.4]
  assign Queue_11_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297341.4]
  assign Queue_11_io_deq_ready = _T_557 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297258.4]
  assign Queue_12_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296480.4]
  assign Queue_12_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296481.4]
  assign Queue_12_io_enq_valid = _T_582 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297343.4]
  assign Queue_12_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297344.4]
  assign Queue_12_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297344.4]
  assign Queue_12_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297344.4]
  assign Queue_12_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297344.4]
  assign Queue_12_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297344.4]
  assign Queue_12_io_deq_ready = _T_586 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297261.4]
  assign Queue_13_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296484.4]
  assign Queue_13_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296485.4]
  assign Queue_13_io_enq_valid = _T_611 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297346.4]
  assign Queue_13_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297347.4]
  assign Queue_13_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297347.4]
  assign Queue_13_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297347.4]
  assign Queue_13_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297347.4]
  assign Queue_13_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297347.4]
  assign Queue_13_io_deq_ready = _T_615 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297264.4]
  assign Queue_14_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296488.4]
  assign Queue_14_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296489.4]
  assign Queue_14_io_enq_valid = _T_640 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297349.4]
  assign Queue_14_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297350.4]
  assign Queue_14_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297350.4]
  assign Queue_14_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297350.4]
  assign Queue_14_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297350.4]
  assign Queue_14_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297350.4]
  assign Queue_14_io_deq_ready = _T_644 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297267.4]
  assign Queue_15_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296492.4]
  assign Queue_15_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296493.4]
  assign Queue_15_io_enq_valid = _T_669 & auto_out_r_valid; // @[Deinterleaver.scala 92:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297352.4]
  assign Queue_15_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297353.4]
  assign Queue_15_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297353.4]
  assign Queue_15_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297353.4]
  assign Queue_15_io_enq_bits_user = auto_out_r_bits_user; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297353.4]
  assign Queue_15_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 93:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297353.4]
  assign Queue_15_io_deq_ready = _T_673 & _T_239; // @[Deinterleaver.scala 86:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297270.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_222 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_224 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_232 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_261 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_290 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_319 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_348 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_377 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_406 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_435 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_464 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_493 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_522 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_551 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_580 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_609 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_638 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_667 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_222 <= 1'h0;
    end else begin
      if (_T_729) begin
        _T_222 <= _T_730;
      end
    end
    _T_224 <= _GEN_1[3:0];
    if (reset) begin
      _T_232 <= 4'h0;
    end else begin
      _T_232 <= _T_246;
    end
    if (reset) begin
      _T_261 <= 4'h0;
    end else begin
      _T_261 <= _T_275;
    end
    if (reset) begin
      _T_290 <= 4'h0;
    end else begin
      _T_290 <= _T_304;
    end
    if (reset) begin
      _T_319 <= 4'h0;
    end else begin
      _T_319 <= _T_333;
    end
    if (reset) begin
      _T_348 <= 4'h0;
    end else begin
      _T_348 <= _T_362;
    end
    if (reset) begin
      _T_377 <= 4'h0;
    end else begin
      _T_377 <= _T_391;
    end
    if (reset) begin
      _T_406 <= 4'h0;
    end else begin
      _T_406 <= _T_420;
    end
    if (reset) begin
      _T_435 <= 4'h0;
    end else begin
      _T_435 <= _T_449;
    end
    if (reset) begin
      _T_464 <= 4'h0;
    end else begin
      _T_464 <= _T_478;
    end
    if (reset) begin
      _T_493 <= 4'h0;
    end else begin
      _T_493 <= _T_507;
    end
    if (reset) begin
      _T_522 <= 4'h0;
    end else begin
      _T_522 <= _T_536;
    end
    if (reset) begin
      _T_551 <= 4'h0;
    end else begin
      _T_551 <= _T_565;
    end
    if (reset) begin
      _T_580 <= 4'h0;
    end else begin
      _T_580 <= _T_594;
    end
    if (reset) begin
      _T_609 <= 4'h0;
    end else begin
      _T_609 <= _T_623;
    end
    if (reset) begin
      _T_638 <= 4'h0;
    end else begin
      _T_638 <= _T_652;
    end
    if (reset) begin
      _T_667 <= 4'h0;
    end else begin
      _T_667 <= _T_681;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_252) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296527.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_252) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296528.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_258) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296537.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_258) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296538.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_281) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296566.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_281) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296567.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_287) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296576.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_287) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296577.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_310) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296605.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_310) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296606.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_316) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296615.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_316) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296616.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_339) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296644.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_339) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296645.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_345) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296654.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_345) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296655.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_368) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296683.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_368) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296684.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_374) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296693.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_374) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296694.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_397) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296722.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_397) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296723.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_403) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296732.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_403) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296733.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_426) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296761.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_426) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296762.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_432) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296771.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_432) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296772.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_455) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296800.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_455) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296801.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_461) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296810.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_461) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296811.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_484) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296839.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_484) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296840.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_490) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296849.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_490) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296850.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_513) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296878.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_513) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296879.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_519) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296888.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_519) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296889.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_542) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296917.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_542) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296918.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_548) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296927.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_548) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296928.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_571) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296956.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_571) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296957.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_577) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296966.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_577) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296967.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296995.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@296996.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_606) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297005.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_606) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297006.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_629) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297034.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_629) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297035.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_635) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297044.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_635) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297045.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_658) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297073.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_658) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297074.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297083.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297084.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_687) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297112.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_687) begin
          $fatal; // @[Deinterleaver.scala 69:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297113.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297122.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693) begin
          $fatal; // @[Deinterleaver.scala 70:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297123.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_62( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297355.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297356.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297357.4]
  output        io_enq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297358.4]
  input         io_enq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297358.4]
  input  [12:0] io_enq_bits, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297358.4]
  input         io_deq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297358.4]
  output        io_deq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297358.4]
  output [12:0] io_deq_bits // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297358.4]
);
  reg [12:0] _T_35 [0:7]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_35__T_58_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
  wire [2:0] _T_35__T_58_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
  wire [12:0] _T_35__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
  wire [2:0] _T_35__T_50_addr; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
  wire  _T_35__T_50_mask; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
  wire  _T_35__T_50_en; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
  reg [2:0] value; // @[Counter.scala 26:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297364.4]
  reg [31:0] _RAND_1;
  reg [2:0] value_1; // @[Counter.scala 26:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297365.4]
  reg [31:0] _RAND_2;
  reg  _T_39; // @[Decoupled.scala 217:35:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297366.4]
  reg [31:0] _RAND_3;
  wire  _T_40; // @[Decoupled.scala 219:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297367.4]
  wire  _T_41; // @[Decoupled.scala 220:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297368.4]
  wire  _T_42; // @[Decoupled.scala 220:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297369.4]
  wire  _T_43; // @[Decoupled.scala 221:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297370.4]
  wire  _T_44; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297371.4]
  wire  _T_47; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297375.4]
  wire [2:0] _T_52; // @[Counter.scala 35:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297384.6]
  wire [2:0] _T_54; // @[Counter.scala 35:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297390.6]
  wire  _T_55; // @[Decoupled.scala 232:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297393.4]
  assign _T_35__T_58_addr = value_1;
  assign _T_35__T_58_data = _T_35[_T_35__T_58_addr]; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
  assign _T_35__T_50_data = io_enq_bits;
  assign _T_35__T_50_addr = value;
  assign _T_35__T_50_mask = 1'h1;
  assign _T_35__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_40 = value == value_1; // @[Decoupled.scala 219:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297367.4]
  assign _T_41 = _T_39 == 1'h0; // @[Decoupled.scala 220:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297368.4]
  assign _T_42 = _T_40 & _T_41; // @[Decoupled.scala 220:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297369.4]
  assign _T_43 = _T_40 & _T_39; // @[Decoupled.scala 221:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297370.4]
  assign _T_44 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297371.4]
  assign _T_47 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297375.4]
  assign _T_52 = value + 3'h1; // @[Counter.scala 35:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297384.6]
  assign _T_54 = value_1 + 3'h1; // @[Counter.scala 35:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297390.6]
  assign _T_55 = _T_44 != _T_47; // @[Decoupled.scala 232:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297393.4]
  assign io_enq_ready = _T_43 == 1'h0; // @[Decoupled.scala 237:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297400.4]
  assign io_deq_valid = _T_42 == 1'h0; // @[Decoupled.scala 236:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297398.4]
  assign io_deq_bits = _T_35__T_58_data; // @[Decoupled.scala 238:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297402.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_35[initvar] = _RAND_0[12:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_39 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35__T_50_en & _T_35__T_50_mask) begin
      _T_35[_T_35__T_50_addr] <= _T_35__T_50_data; // @[Decoupled.scala 214:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@297363.4]
    end
    if (reset) begin
      value <= 3'h0;
    end else begin
      if (_T_44) begin
        value <= _T_52;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (_T_47) begin
        value_1 <= _T_54;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_55) begin
        _T_39 <= _T_44;
      end
    end
  end
endmodule
module AXI4UserYanker( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299115.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299116.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299117.4]
  output        auto_in_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_in_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [3:0]  auto_in_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [31:0] auto_in_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_in_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [12:0] auto_in_aw_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_in_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_in_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [63:0] auto_in_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [7:0]  auto_in_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_in_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_in_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_in_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [3:0]  auto_in_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [1:0]  auto_in_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [12:0] auto_in_b_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_in_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_in_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [3:0]  auto_in_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [31:0] auto_in_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_in_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [12:0] auto_in_ar_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_in_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_in_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [3:0]  auto_in_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [63:0] auto_in_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [1:0]  auto_in_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [12:0] auto_in_r_bits_user, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_in_r_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_out_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_out_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [3:0]  auto_out_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [31:0] auto_out_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [7:0]  auto_out_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [2:0]  auto_out_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_out_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_out_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_out_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [63:0] auto_out_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [7:0]  auto_out_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_out_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_out_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_out_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [3:0]  auto_out_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_out_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_out_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [3:0]  auto_out_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [31:0] auto_out_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [7:0]  auto_out_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [2:0]  auto_out_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_out_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  output        auto_out_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_out_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [3:0]  auto_out_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [63:0] auto_out_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
  input         auto_out_r_bits_last // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299118.4]
);
  wire  Queue_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
  wire  Queue_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
  wire  Queue_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
  wire  Queue_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
  wire [12:0] Queue_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
  wire  Queue_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
  wire  Queue_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
  wire [12:0] Queue_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
  wire  Queue_1_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
  wire  Queue_1_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
  wire  Queue_1_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
  wire  Queue_1_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
  wire [12:0] Queue_1_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
  wire  Queue_1_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
  wire  Queue_1_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
  wire [12:0] Queue_1_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
  wire  Queue_2_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
  wire  Queue_2_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
  wire  Queue_2_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
  wire  Queue_2_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
  wire [12:0] Queue_2_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
  wire  Queue_2_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
  wire  Queue_2_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
  wire [12:0] Queue_2_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
  wire  Queue_3_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
  wire  Queue_3_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
  wire  Queue_3_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
  wire  Queue_3_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
  wire [12:0] Queue_3_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
  wire  Queue_3_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
  wire  Queue_3_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
  wire [12:0] Queue_3_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
  wire  Queue_4_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
  wire  Queue_4_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
  wire  Queue_4_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
  wire  Queue_4_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
  wire [12:0] Queue_4_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
  wire  Queue_4_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
  wire  Queue_4_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
  wire [12:0] Queue_4_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
  wire  Queue_5_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
  wire  Queue_5_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
  wire  Queue_5_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
  wire  Queue_5_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
  wire [12:0] Queue_5_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
  wire  Queue_5_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
  wire  Queue_5_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
  wire [12:0] Queue_5_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
  wire  Queue_6_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
  wire  Queue_6_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
  wire  Queue_6_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
  wire  Queue_6_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
  wire [12:0] Queue_6_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
  wire  Queue_6_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
  wire  Queue_6_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
  wire [12:0] Queue_6_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
  wire  Queue_7_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
  wire  Queue_7_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
  wire  Queue_7_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
  wire  Queue_7_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
  wire [12:0] Queue_7_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
  wire  Queue_7_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
  wire  Queue_7_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
  wire [12:0] Queue_7_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
  wire  Queue_8_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
  wire  Queue_8_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
  wire  Queue_8_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
  wire  Queue_8_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
  wire [12:0] Queue_8_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
  wire  Queue_8_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
  wire  Queue_8_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
  wire [12:0] Queue_8_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
  wire  Queue_9_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
  wire  Queue_9_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
  wire  Queue_9_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
  wire  Queue_9_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
  wire [12:0] Queue_9_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
  wire  Queue_9_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
  wire  Queue_9_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
  wire [12:0] Queue_9_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
  wire  Queue_10_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
  wire  Queue_10_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
  wire  Queue_10_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
  wire  Queue_10_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
  wire [12:0] Queue_10_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
  wire  Queue_10_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
  wire  Queue_10_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
  wire [12:0] Queue_10_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
  wire  Queue_11_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
  wire  Queue_11_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
  wire  Queue_11_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
  wire  Queue_11_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
  wire [12:0] Queue_11_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
  wire  Queue_11_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
  wire  Queue_11_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
  wire [12:0] Queue_11_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
  wire  Queue_12_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
  wire  Queue_12_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
  wire  Queue_12_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
  wire  Queue_12_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
  wire [12:0] Queue_12_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
  wire  Queue_12_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
  wire  Queue_12_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
  wire [12:0] Queue_12_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
  wire  Queue_13_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
  wire  Queue_13_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
  wire  Queue_13_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
  wire  Queue_13_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
  wire [12:0] Queue_13_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
  wire  Queue_13_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
  wire  Queue_13_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
  wire [12:0] Queue_13_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
  wire  Queue_14_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
  wire  Queue_14_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
  wire  Queue_14_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
  wire  Queue_14_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
  wire [12:0] Queue_14_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
  wire  Queue_14_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
  wire  Queue_14_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
  wire [12:0] Queue_14_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
  wire  Queue_15_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
  wire  Queue_15_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
  wire  Queue_15_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
  wire  Queue_15_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
  wire [12:0] Queue_15_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
  wire  Queue_15_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
  wire  Queue_15_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
  wire [12:0] Queue_15_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
  wire  Queue_16_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
  wire  Queue_16_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
  wire  Queue_16_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
  wire  Queue_16_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
  wire [12:0] Queue_16_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
  wire  Queue_16_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
  wire  Queue_16_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
  wire [12:0] Queue_16_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
  wire  Queue_17_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
  wire  Queue_17_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
  wire  Queue_17_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
  wire  Queue_17_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
  wire [12:0] Queue_17_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
  wire  Queue_17_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
  wire  Queue_17_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
  wire [12:0] Queue_17_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
  wire  Queue_18_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
  wire  Queue_18_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
  wire  Queue_18_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
  wire  Queue_18_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
  wire [12:0] Queue_18_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
  wire  Queue_18_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
  wire  Queue_18_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
  wire [12:0] Queue_18_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
  wire  Queue_19_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
  wire  Queue_19_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
  wire  Queue_19_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
  wire  Queue_19_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
  wire [12:0] Queue_19_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
  wire  Queue_19_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
  wire  Queue_19_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
  wire [12:0] Queue_19_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
  wire  Queue_20_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
  wire  Queue_20_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
  wire  Queue_20_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
  wire  Queue_20_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
  wire [12:0] Queue_20_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
  wire  Queue_20_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
  wire  Queue_20_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
  wire [12:0] Queue_20_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
  wire  Queue_21_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
  wire  Queue_21_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
  wire  Queue_21_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
  wire  Queue_21_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
  wire [12:0] Queue_21_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
  wire  Queue_21_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
  wire  Queue_21_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
  wire [12:0] Queue_21_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
  wire  Queue_22_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
  wire  Queue_22_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
  wire  Queue_22_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
  wire  Queue_22_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
  wire [12:0] Queue_22_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
  wire  Queue_22_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
  wire  Queue_22_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
  wire [12:0] Queue_22_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
  wire  Queue_23_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
  wire  Queue_23_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
  wire  Queue_23_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
  wire  Queue_23_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
  wire [12:0] Queue_23_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
  wire  Queue_23_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
  wire  Queue_23_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
  wire [12:0] Queue_23_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
  wire  Queue_24_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
  wire  Queue_24_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
  wire  Queue_24_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
  wire  Queue_24_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
  wire [12:0] Queue_24_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
  wire  Queue_24_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
  wire  Queue_24_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
  wire [12:0] Queue_24_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
  wire  Queue_25_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
  wire  Queue_25_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
  wire  Queue_25_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
  wire  Queue_25_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
  wire [12:0] Queue_25_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
  wire  Queue_25_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
  wire  Queue_25_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
  wire [12:0] Queue_25_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
  wire  Queue_26_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
  wire  Queue_26_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
  wire  Queue_26_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
  wire  Queue_26_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
  wire [12:0] Queue_26_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
  wire  Queue_26_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
  wire  Queue_26_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
  wire [12:0] Queue_26_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
  wire  Queue_27_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
  wire  Queue_27_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
  wire  Queue_27_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
  wire  Queue_27_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
  wire [12:0] Queue_27_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
  wire  Queue_27_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
  wire  Queue_27_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
  wire [12:0] Queue_27_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
  wire  Queue_28_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
  wire  Queue_28_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
  wire  Queue_28_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
  wire  Queue_28_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
  wire [12:0] Queue_28_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
  wire  Queue_28_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
  wire  Queue_28_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
  wire [12:0] Queue_28_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
  wire  Queue_29_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
  wire  Queue_29_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
  wire  Queue_29_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
  wire  Queue_29_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
  wire [12:0] Queue_29_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
  wire  Queue_29_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
  wire  Queue_29_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
  wire [12:0] Queue_29_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
  wire  Queue_30_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
  wire  Queue_30_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
  wire  Queue_30_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
  wire  Queue_30_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
  wire [12:0] Queue_30_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
  wire  Queue_30_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
  wire  Queue_30_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
  wire [12:0] Queue_30_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
  wire  Queue_31_clock; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
  wire  Queue_31_reset; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
  wire  Queue_31_io_enq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
  wire  Queue_31_io_enq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
  wire [12:0] Queue_31_io_enq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
  wire  Queue_31_io_deq_ready; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
  wire  Queue_31_io_deq_valid; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
  wire [12:0] Queue_31_io_deq_bits; // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
  wire  _T_224_0; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299259.4]
  wire  _T_224_1; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299260.4]
  wire  _GEN_1; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_2; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299261.4]
  wire  _GEN_2; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_3; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299262.4]
  wire  _GEN_3; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_4; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299263.4]
  wire  _GEN_4; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_5; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299264.4]
  wire  _GEN_5; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_6; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299265.4]
  wire  _GEN_6; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_7; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299266.4]
  wire  _GEN_7; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_8; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299267.4]
  wire  _GEN_8; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_9; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299268.4]
  wire  _GEN_9; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_10; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299269.4]
  wire  _GEN_10; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_11; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299270.4]
  wire  _GEN_11; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_12; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299271.4]
  wire  _GEN_12; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_13; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299272.4]
  wire  _GEN_13; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_14; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299273.4]
  wire  _GEN_14; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_224_15; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299274.4]
  wire  _GEN_15; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  wire  _T_292; // @[UserYanker.scala 54:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299316.4]
  wire  _T_249_0; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299282.4]
  wire  _T_249_1; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299283.4]
  wire  _GEN_17; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_2; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299284.4]
  wire  _GEN_18; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_3; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299285.4]
  wire  _GEN_19; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_4; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299286.4]
  wire  _GEN_20; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_5; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299287.4]
  wire  _GEN_21; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_6; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299288.4]
  wire  _GEN_22; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_7; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299289.4]
  wire  _GEN_23; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_8; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299290.4]
  wire  _GEN_24; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_9; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299291.4]
  wire  _GEN_25; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_10; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299292.4]
  wire  _GEN_26; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_11; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299293.4]
  wire  _GEN_27; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_12; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299294.4]
  wire  _GEN_28; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_13; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299295.4]
  wire  _GEN_29; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_14; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299296.4]
  wire  _GEN_30; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_249_15; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299297.4]
  wire  _GEN_31; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_293; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  wire  _T_295; // @[UserYanker.scala 54:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299319.4]
  wire  _T_296; // @[UserYanker.scala 54:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299320.4]
  wire [12:0] _T_272_0; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299300.4]
  wire [12:0] _T_272_1; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299301.4]
  wire [12:0] _GEN_33; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_2; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299302.4]
  wire [12:0] _GEN_34; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_3; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299303.4]
  wire [12:0] _GEN_35; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_4; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299304.4]
  wire [12:0] _GEN_36; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_5; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299305.4]
  wire [12:0] _GEN_37; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_6; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299306.4]
  wire [12:0] _GEN_38; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_7; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299307.4]
  wire [12:0] _GEN_39; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_8; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299308.4]
  wire [12:0] _GEN_40; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_9; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299309.4]
  wire [12:0] _GEN_41; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_10; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299310.4]
  wire [12:0] _GEN_42; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_11; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299311.4]
  wire [12:0] _GEN_43; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_12; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299312.4]
  wire [12:0] _GEN_44; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_13; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299313.4]
  wire [12:0] _GEN_45; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_14; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299314.4]
  wire [12:0] _GEN_46; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  wire [12:0] _T_272_15; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299315.4]
  wire [15:0] _T_298; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299328.4]
  wire  _T_300; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299330.4]
  wire  _T_301; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299331.4]
  wire  _T_302; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299332.4]
  wire  _T_303; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299333.4]
  wire  _T_304; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299334.4]
  wire  _T_305; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299335.4]
  wire  _T_306; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299336.4]
  wire  _T_307; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299337.4]
  wire  _T_308; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299338.4]
  wire  _T_309; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299339.4]
  wire  _T_310; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299340.4]
  wire  _T_311; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299341.4]
  wire  _T_312; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299342.4]
  wire  _T_313; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299343.4]
  wire  _T_314; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299344.4]
  wire  _T_315; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299345.4]
  wire [15:0] _T_317; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299347.4]
  wire  _T_319; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299349.4]
  wire  _T_320; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299350.4]
  wire  _T_321; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299351.4]
  wire  _T_322; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299352.4]
  wire  _T_323; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299353.4]
  wire  _T_324; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299354.4]
  wire  _T_325; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299355.4]
  wire  _T_326; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299356.4]
  wire  _T_327; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299357.4]
  wire  _T_328; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299358.4]
  wire  _T_329; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299359.4]
  wire  _T_330; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299360.4]
  wire  _T_331; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299361.4]
  wire  _T_332; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299362.4]
  wire  _T_333; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299363.4]
  wire  _T_334; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299364.4]
  wire  _T_335; // @[UserYanker.scala 61:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299365.4]
  wire  _T_336; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299366.4]
  wire  _T_338; // @[UserYanker.scala 62:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299369.4]
  wire  _T_341; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299374.4]
  wire  _T_346; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299382.4]
  wire  _T_351; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299390.4]
  wire  _T_356; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299398.4]
  wire  _T_361; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299406.4]
  wire  _T_366; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299414.4]
  wire  _T_371; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299422.4]
  wire  _T_376; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299430.4]
  wire  _T_381; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299438.4]
  wire  _T_386; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299446.4]
  wire  _T_391; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299454.4]
  wire  _T_396; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299462.4]
  wire  _T_401; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299470.4]
  wire  _T_406; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299478.4]
  wire  _T_411; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299486.4]
  wire  _T_418_0; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299495.4]
  wire  _T_418_1; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299496.4]
  wire  _GEN_49; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_2; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299497.4]
  wire  _GEN_50; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_3; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299498.4]
  wire  _GEN_51; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_4; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299499.4]
  wire  _GEN_52; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_5; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299500.4]
  wire  _GEN_53; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_6; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299501.4]
  wire  _GEN_54; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_7; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299502.4]
  wire  _GEN_55; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_8; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299503.4]
  wire  _GEN_56; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_9; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299504.4]
  wire  _GEN_57; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_10; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299505.4]
  wire  _GEN_58; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_11; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299506.4]
  wire  _GEN_59; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_12; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299507.4]
  wire  _GEN_60; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_13; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299508.4]
  wire  _GEN_61; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_14; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299509.4]
  wire  _GEN_62; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_418_15; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299510.4]
  wire  _GEN_63; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  wire  _T_486; // @[UserYanker.scala 75:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299552.4]
  wire  _T_443_0; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299518.4]
  wire  _T_443_1; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299519.4]
  wire  _GEN_65; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_2; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299520.4]
  wire  _GEN_66; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_3; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299521.4]
  wire  _GEN_67; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_4; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299522.4]
  wire  _GEN_68; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_5; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299523.4]
  wire  _GEN_69; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_6; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299524.4]
  wire  _GEN_70; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_7; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299525.4]
  wire  _GEN_71; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_8; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299526.4]
  wire  _GEN_72; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_9; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299527.4]
  wire  _GEN_73; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_10; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299528.4]
  wire  _GEN_74; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_11; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299529.4]
  wire  _GEN_75; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_12; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299530.4]
  wire  _GEN_76; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_13; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299531.4]
  wire  _GEN_77; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_14; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299532.4]
  wire  _GEN_78; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_443_15; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299533.4]
  wire  _GEN_79; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_487; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  wire  _T_489; // @[UserYanker.scala 75:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299555.4]
  wire  _T_490; // @[UserYanker.scala 75:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299556.4]
  wire [12:0] _T_466_0; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299536.4]
  wire [12:0] _T_466_1; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299537.4]
  wire [12:0] _GEN_81; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_2; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299538.4]
  wire [12:0] _GEN_82; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_3; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299539.4]
  wire [12:0] _GEN_83; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_4; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299540.4]
  wire [12:0] _GEN_84; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_5; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299541.4]
  wire [12:0] _GEN_85; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_6; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299542.4]
  wire [12:0] _GEN_86; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_7; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299543.4]
  wire [12:0] _GEN_87; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_8; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299544.4]
  wire [12:0] _GEN_88; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_9; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299545.4]
  wire [12:0] _GEN_89; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_10; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299546.4]
  wire [12:0] _GEN_90; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_11; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299547.4]
  wire [12:0] _GEN_91; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_12; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299548.4]
  wire [12:0] _GEN_92; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_13; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299549.4]
  wire [12:0] _GEN_93; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_14; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299550.4]
  wire [12:0] _GEN_94; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  wire [12:0] _T_466_15; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299551.4]
  wire [15:0] _T_492; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299564.4]
  wire  _T_494; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299566.4]
  wire  _T_495; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299567.4]
  wire  _T_496; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299568.4]
  wire  _T_497; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299569.4]
  wire  _T_498; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299570.4]
  wire  _T_499; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299571.4]
  wire  _T_500; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299572.4]
  wire  _T_501; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299573.4]
  wire  _T_502; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299574.4]
  wire  _T_503; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299575.4]
  wire  _T_504; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299576.4]
  wire  _T_505; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299577.4]
  wire  _T_506; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299578.4]
  wire  _T_507; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299579.4]
  wire  _T_508; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299580.4]
  wire  _T_509; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299581.4]
  wire [15:0] _T_511; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299583.4]
  wire  _T_513; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299585.4]
  wire  _T_514; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299586.4]
  wire  _T_515; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299587.4]
  wire  _T_516; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299588.4]
  wire  _T_517; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299589.4]
  wire  _T_518; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299590.4]
  wire  _T_519; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299591.4]
  wire  _T_520; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299592.4]
  wire  _T_521; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299593.4]
  wire  _T_522; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299594.4]
  wire  _T_523; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299595.4]
  wire  _T_524; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299596.4]
  wire  _T_525; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299597.4]
  wire  _T_526; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299598.4]
  wire  _T_527; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299599.4]
  wire  _T_528; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299600.4]
  wire  _T_529; // @[UserYanker.scala 82:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299601.4]
  wire  _T_531; // @[UserYanker.scala 83:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299604.4]
  Queue_62 Queue ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299129.4]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  Queue_62 Queue_1 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299133.4]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  Queue_62 Queue_2 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299137.4]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  Queue_62 Queue_3 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299141.4]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  Queue_62 Queue_4 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299145.4]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits(Queue_4_io_enq_bits),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits(Queue_4_io_deq_bits)
  );
  Queue_62 Queue_5 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299149.4]
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits(Queue_5_io_enq_bits),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits(Queue_5_io_deq_bits)
  );
  Queue_62 Queue_6 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299153.4]
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits(Queue_6_io_enq_bits),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits(Queue_6_io_deq_bits)
  );
  Queue_62 Queue_7 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299157.4]
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits(Queue_7_io_enq_bits),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits(Queue_7_io_deq_bits)
  );
  Queue_62 Queue_8 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299161.4]
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits(Queue_8_io_enq_bits),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits(Queue_8_io_deq_bits)
  );
  Queue_62 Queue_9 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299165.4]
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits(Queue_9_io_enq_bits),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits(Queue_9_io_deq_bits)
  );
  Queue_62 Queue_10 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299169.4]
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits(Queue_10_io_enq_bits),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits(Queue_10_io_deq_bits)
  );
  Queue_62 Queue_11 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299173.4]
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits(Queue_11_io_enq_bits),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits(Queue_11_io_deq_bits)
  );
  Queue_62 Queue_12 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299177.4]
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits(Queue_12_io_enq_bits),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits(Queue_12_io_deq_bits)
  );
  Queue_62 Queue_13 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299181.4]
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits(Queue_13_io_enq_bits),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits(Queue_13_io_deq_bits)
  );
  Queue_62 Queue_14 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299185.4]
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits(Queue_14_io_enq_bits),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits(Queue_14_io_deq_bits)
  );
  Queue_62 Queue_15 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299189.4]
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits(Queue_15_io_enq_bits),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits(Queue_15_io_deq_bits)
  );
  Queue_62 Queue_16 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299193.4]
    .clock(Queue_16_clock),
    .reset(Queue_16_reset),
    .io_enq_ready(Queue_16_io_enq_ready),
    .io_enq_valid(Queue_16_io_enq_valid),
    .io_enq_bits(Queue_16_io_enq_bits),
    .io_deq_ready(Queue_16_io_deq_ready),
    .io_deq_valid(Queue_16_io_deq_valid),
    .io_deq_bits(Queue_16_io_deq_bits)
  );
  Queue_62 Queue_17 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299197.4]
    .clock(Queue_17_clock),
    .reset(Queue_17_reset),
    .io_enq_ready(Queue_17_io_enq_ready),
    .io_enq_valid(Queue_17_io_enq_valid),
    .io_enq_bits(Queue_17_io_enq_bits),
    .io_deq_ready(Queue_17_io_deq_ready),
    .io_deq_valid(Queue_17_io_deq_valid),
    .io_deq_bits(Queue_17_io_deq_bits)
  );
  Queue_62 Queue_18 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299201.4]
    .clock(Queue_18_clock),
    .reset(Queue_18_reset),
    .io_enq_ready(Queue_18_io_enq_ready),
    .io_enq_valid(Queue_18_io_enq_valid),
    .io_enq_bits(Queue_18_io_enq_bits),
    .io_deq_ready(Queue_18_io_deq_ready),
    .io_deq_valid(Queue_18_io_deq_valid),
    .io_deq_bits(Queue_18_io_deq_bits)
  );
  Queue_62 Queue_19 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299205.4]
    .clock(Queue_19_clock),
    .reset(Queue_19_reset),
    .io_enq_ready(Queue_19_io_enq_ready),
    .io_enq_valid(Queue_19_io_enq_valid),
    .io_enq_bits(Queue_19_io_enq_bits),
    .io_deq_ready(Queue_19_io_deq_ready),
    .io_deq_valid(Queue_19_io_deq_valid),
    .io_deq_bits(Queue_19_io_deq_bits)
  );
  Queue_62 Queue_20 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299209.4]
    .clock(Queue_20_clock),
    .reset(Queue_20_reset),
    .io_enq_ready(Queue_20_io_enq_ready),
    .io_enq_valid(Queue_20_io_enq_valid),
    .io_enq_bits(Queue_20_io_enq_bits),
    .io_deq_ready(Queue_20_io_deq_ready),
    .io_deq_valid(Queue_20_io_deq_valid),
    .io_deq_bits(Queue_20_io_deq_bits)
  );
  Queue_62 Queue_21 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299213.4]
    .clock(Queue_21_clock),
    .reset(Queue_21_reset),
    .io_enq_ready(Queue_21_io_enq_ready),
    .io_enq_valid(Queue_21_io_enq_valid),
    .io_enq_bits(Queue_21_io_enq_bits),
    .io_deq_ready(Queue_21_io_deq_ready),
    .io_deq_valid(Queue_21_io_deq_valid),
    .io_deq_bits(Queue_21_io_deq_bits)
  );
  Queue_62 Queue_22 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299217.4]
    .clock(Queue_22_clock),
    .reset(Queue_22_reset),
    .io_enq_ready(Queue_22_io_enq_ready),
    .io_enq_valid(Queue_22_io_enq_valid),
    .io_enq_bits(Queue_22_io_enq_bits),
    .io_deq_ready(Queue_22_io_deq_ready),
    .io_deq_valid(Queue_22_io_deq_valid),
    .io_deq_bits(Queue_22_io_deq_bits)
  );
  Queue_62 Queue_23 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299221.4]
    .clock(Queue_23_clock),
    .reset(Queue_23_reset),
    .io_enq_ready(Queue_23_io_enq_ready),
    .io_enq_valid(Queue_23_io_enq_valid),
    .io_enq_bits(Queue_23_io_enq_bits),
    .io_deq_ready(Queue_23_io_deq_ready),
    .io_deq_valid(Queue_23_io_deq_valid),
    .io_deq_bits(Queue_23_io_deq_bits)
  );
  Queue_62 Queue_24 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299225.4]
    .clock(Queue_24_clock),
    .reset(Queue_24_reset),
    .io_enq_ready(Queue_24_io_enq_ready),
    .io_enq_valid(Queue_24_io_enq_valid),
    .io_enq_bits(Queue_24_io_enq_bits),
    .io_deq_ready(Queue_24_io_deq_ready),
    .io_deq_valid(Queue_24_io_deq_valid),
    .io_deq_bits(Queue_24_io_deq_bits)
  );
  Queue_62 Queue_25 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299229.4]
    .clock(Queue_25_clock),
    .reset(Queue_25_reset),
    .io_enq_ready(Queue_25_io_enq_ready),
    .io_enq_valid(Queue_25_io_enq_valid),
    .io_enq_bits(Queue_25_io_enq_bits),
    .io_deq_ready(Queue_25_io_deq_ready),
    .io_deq_valid(Queue_25_io_deq_valid),
    .io_deq_bits(Queue_25_io_deq_bits)
  );
  Queue_62 Queue_26 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299233.4]
    .clock(Queue_26_clock),
    .reset(Queue_26_reset),
    .io_enq_ready(Queue_26_io_enq_ready),
    .io_enq_valid(Queue_26_io_enq_valid),
    .io_enq_bits(Queue_26_io_enq_bits),
    .io_deq_ready(Queue_26_io_deq_ready),
    .io_deq_valid(Queue_26_io_deq_valid),
    .io_deq_bits(Queue_26_io_deq_bits)
  );
  Queue_62 Queue_27 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299237.4]
    .clock(Queue_27_clock),
    .reset(Queue_27_reset),
    .io_enq_ready(Queue_27_io_enq_ready),
    .io_enq_valid(Queue_27_io_enq_valid),
    .io_enq_bits(Queue_27_io_enq_bits),
    .io_deq_ready(Queue_27_io_deq_ready),
    .io_deq_valid(Queue_27_io_deq_valid),
    .io_deq_bits(Queue_27_io_deq_bits)
  );
  Queue_62 Queue_28 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299241.4]
    .clock(Queue_28_clock),
    .reset(Queue_28_reset),
    .io_enq_ready(Queue_28_io_enq_ready),
    .io_enq_valid(Queue_28_io_enq_valid),
    .io_enq_bits(Queue_28_io_enq_bits),
    .io_deq_ready(Queue_28_io_deq_ready),
    .io_deq_valid(Queue_28_io_deq_valid),
    .io_deq_bits(Queue_28_io_deq_bits)
  );
  Queue_62 Queue_29 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299245.4]
    .clock(Queue_29_clock),
    .reset(Queue_29_reset),
    .io_enq_ready(Queue_29_io_enq_ready),
    .io_enq_valid(Queue_29_io_enq_valid),
    .io_enq_bits(Queue_29_io_enq_bits),
    .io_deq_ready(Queue_29_io_deq_ready),
    .io_deq_valid(Queue_29_io_deq_valid),
    .io_deq_bits(Queue_29_io_deq_bits)
  );
  Queue_62 Queue_30 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299249.4]
    .clock(Queue_30_clock),
    .reset(Queue_30_reset),
    .io_enq_ready(Queue_30_io_enq_ready),
    .io_enq_valid(Queue_30_io_enq_valid),
    .io_enq_bits(Queue_30_io_enq_bits),
    .io_deq_ready(Queue_30_io_deq_ready),
    .io_deq_valid(Queue_30_io_deq_valid),
    .io_deq_bits(Queue_30_io_deq_bits)
  );
  Queue_62 Queue_31 ( // @[UserYanker.scala 38:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299253.4]
    .clock(Queue_31_clock),
    .reset(Queue_31_reset),
    .io_enq_ready(Queue_31_io_enq_ready),
    .io_enq_valid(Queue_31_io_enq_valid),
    .io_enq_bits(Queue_31_io_enq_bits),
    .io_deq_ready(Queue_31_io_deq_ready),
    .io_deq_valid(Queue_31_io_deq_valid),
    .io_deq_bits(Queue_31_io_deq_bits)
  );
  assign _T_224_0 = Queue_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299259.4]
  assign _T_224_1 = Queue_1_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299260.4]
  assign _GEN_1 = 4'h1 == auto_in_ar_bits_id ? _T_224_1 : _T_224_0; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_2 = Queue_2_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299261.4]
  assign _GEN_2 = 4'h2 == auto_in_ar_bits_id ? _T_224_2 : _GEN_1; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_3 = Queue_3_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299262.4]
  assign _GEN_3 = 4'h3 == auto_in_ar_bits_id ? _T_224_3 : _GEN_2; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_4 = Queue_4_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299263.4]
  assign _GEN_4 = 4'h4 == auto_in_ar_bits_id ? _T_224_4 : _GEN_3; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_5 = Queue_5_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299264.4]
  assign _GEN_5 = 4'h5 == auto_in_ar_bits_id ? _T_224_5 : _GEN_4; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_6 = Queue_6_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299265.4]
  assign _GEN_6 = 4'h6 == auto_in_ar_bits_id ? _T_224_6 : _GEN_5; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_7 = Queue_7_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299266.4]
  assign _GEN_7 = 4'h7 == auto_in_ar_bits_id ? _T_224_7 : _GEN_6; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_8 = Queue_8_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299267.4]
  assign _GEN_8 = 4'h8 == auto_in_ar_bits_id ? _T_224_8 : _GEN_7; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_9 = Queue_9_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299268.4]
  assign _GEN_9 = 4'h9 == auto_in_ar_bits_id ? _T_224_9 : _GEN_8; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_10 = Queue_10_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299269.4]
  assign _GEN_10 = 4'ha == auto_in_ar_bits_id ? _T_224_10 : _GEN_9; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_11 = Queue_11_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299270.4]
  assign _GEN_11 = 4'hb == auto_in_ar_bits_id ? _T_224_11 : _GEN_10; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_12 = Queue_12_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299271.4]
  assign _GEN_12 = 4'hc == auto_in_ar_bits_id ? _T_224_12 : _GEN_11; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_13 = Queue_13_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299272.4]
  assign _GEN_13 = 4'hd == auto_in_ar_bits_id ? _T_224_13 : _GEN_12; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_14 = Queue_14_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299273.4]
  assign _GEN_14 = 4'he == auto_in_ar_bits_id ? _T_224_14 : _GEN_13; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_224_15 = Queue_15_io_enq_ready; // @[UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299257.4 UserYanker.scala 46:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299274.4]
  assign _GEN_15 = 4'hf == auto_in_ar_bits_id ? _T_224_15 : _GEN_14; // @[UserYanker.scala 47:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299275.4]
  assign _T_292 = auto_out_r_valid == 1'h0; // @[UserYanker.scala 54:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299316.4]
  assign _T_249_0 = Queue_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299282.4]
  assign _T_249_1 = Queue_1_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299283.4]
  assign _GEN_17 = 4'h1 == auto_out_r_bits_id ? _T_249_1 : _T_249_0; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_2 = Queue_2_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299284.4]
  assign _GEN_18 = 4'h2 == auto_out_r_bits_id ? _T_249_2 : _GEN_17; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_3 = Queue_3_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299285.4]
  assign _GEN_19 = 4'h3 == auto_out_r_bits_id ? _T_249_3 : _GEN_18; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_4 = Queue_4_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299286.4]
  assign _GEN_20 = 4'h4 == auto_out_r_bits_id ? _T_249_4 : _GEN_19; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_5 = Queue_5_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299287.4]
  assign _GEN_21 = 4'h5 == auto_out_r_bits_id ? _T_249_5 : _GEN_20; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_6 = Queue_6_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299288.4]
  assign _GEN_22 = 4'h6 == auto_out_r_bits_id ? _T_249_6 : _GEN_21; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_7 = Queue_7_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299289.4]
  assign _GEN_23 = 4'h7 == auto_out_r_bits_id ? _T_249_7 : _GEN_22; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_8 = Queue_8_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299290.4]
  assign _GEN_24 = 4'h8 == auto_out_r_bits_id ? _T_249_8 : _GEN_23; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_9 = Queue_9_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299291.4]
  assign _GEN_25 = 4'h9 == auto_out_r_bits_id ? _T_249_9 : _GEN_24; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_10 = Queue_10_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299292.4]
  assign _GEN_26 = 4'ha == auto_out_r_bits_id ? _T_249_10 : _GEN_25; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_11 = Queue_11_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299293.4]
  assign _GEN_27 = 4'hb == auto_out_r_bits_id ? _T_249_11 : _GEN_26; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_12 = Queue_12_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299294.4]
  assign _GEN_28 = 4'hc == auto_out_r_bits_id ? _T_249_12 : _GEN_27; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_13 = Queue_13_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299295.4]
  assign _GEN_29 = 4'hd == auto_out_r_bits_id ? _T_249_13 : _GEN_28; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_14 = Queue_14_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299296.4]
  assign _GEN_30 = 4'he == auto_out_r_bits_id ? _T_249_14 : _GEN_29; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_249_15 = Queue_15_io_deq_valid; // @[UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299280.4 UserYanker.scala 52:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299297.4]
  assign _GEN_31 = 4'hf == auto_out_r_bits_id ? _T_249_15 : _GEN_30; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_293 = _T_292 | _GEN_31; // @[UserYanker.scala 54:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299317.4]
  assign _T_295 = _T_293 | reset; // @[UserYanker.scala 54:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299319.4]
  assign _T_296 = _T_295 == 1'h0; // @[UserYanker.scala 54:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299320.4]
  assign _T_272_0 = Queue_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299300.4]
  assign _T_272_1 = Queue_1_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299301.4]
  assign _GEN_33 = 4'h1 == auto_out_r_bits_id ? _T_272_1 : _T_272_0; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_2 = Queue_2_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299302.4]
  assign _GEN_34 = 4'h2 == auto_out_r_bits_id ? _T_272_2 : _GEN_33; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_3 = Queue_3_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299303.4]
  assign _GEN_35 = 4'h3 == auto_out_r_bits_id ? _T_272_3 : _GEN_34; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_4 = Queue_4_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299304.4]
  assign _GEN_36 = 4'h4 == auto_out_r_bits_id ? _T_272_4 : _GEN_35; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_5 = Queue_5_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299305.4]
  assign _GEN_37 = 4'h5 == auto_out_r_bits_id ? _T_272_5 : _GEN_36; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_6 = Queue_6_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299306.4]
  assign _GEN_38 = 4'h6 == auto_out_r_bits_id ? _T_272_6 : _GEN_37; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_7 = Queue_7_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299307.4]
  assign _GEN_39 = 4'h7 == auto_out_r_bits_id ? _T_272_7 : _GEN_38; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_8 = Queue_8_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299308.4]
  assign _GEN_40 = 4'h8 == auto_out_r_bits_id ? _T_272_8 : _GEN_39; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_9 = Queue_9_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299309.4]
  assign _GEN_41 = 4'h9 == auto_out_r_bits_id ? _T_272_9 : _GEN_40; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_10 = Queue_10_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299310.4]
  assign _GEN_42 = 4'ha == auto_out_r_bits_id ? _T_272_10 : _GEN_41; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_11 = Queue_11_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299311.4]
  assign _GEN_43 = 4'hb == auto_out_r_bits_id ? _T_272_11 : _GEN_42; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_12 = Queue_12_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299312.4]
  assign _GEN_44 = 4'hc == auto_out_r_bits_id ? _T_272_12 : _GEN_43; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_13 = Queue_13_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299313.4]
  assign _GEN_45 = 4'hd == auto_out_r_bits_id ? _T_272_13 : _GEN_44; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_14 = Queue_14_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299314.4]
  assign _GEN_46 = 4'he == auto_out_r_bits_id ? _T_272_14 : _GEN_45; // @[UserYanker.scala 56:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299326.4]
  assign _T_272_15 = Queue_15_io_deq_bits; // @[UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299298.4 UserYanker.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299315.4]
  assign _T_298 = 16'h1 << auto_in_ar_bits_id; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299328.4]
  assign _T_300 = _T_298[0]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299330.4]
  assign _T_301 = _T_298[1]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299331.4]
  assign _T_302 = _T_298[2]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299332.4]
  assign _T_303 = _T_298[3]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299333.4]
  assign _T_304 = _T_298[4]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299334.4]
  assign _T_305 = _T_298[5]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299335.4]
  assign _T_306 = _T_298[6]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299336.4]
  assign _T_307 = _T_298[7]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299337.4]
  assign _T_308 = _T_298[8]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299338.4]
  assign _T_309 = _T_298[9]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299339.4]
  assign _T_310 = _T_298[10]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299340.4]
  assign _T_311 = _T_298[11]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299341.4]
  assign _T_312 = _T_298[12]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299342.4]
  assign _T_313 = _T_298[13]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299343.4]
  assign _T_314 = _T_298[14]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299344.4]
  assign _T_315 = _T_298[15]; // @[UserYanker.scala 58:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299345.4]
  assign _T_317 = 16'h1 << auto_out_r_bits_id; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299347.4]
  assign _T_319 = _T_317[0]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299349.4]
  assign _T_320 = _T_317[1]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299350.4]
  assign _T_321 = _T_317[2]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299351.4]
  assign _T_322 = _T_317[3]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299352.4]
  assign _T_323 = _T_317[4]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299353.4]
  assign _T_324 = _T_317[5]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299354.4]
  assign _T_325 = _T_317[6]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299355.4]
  assign _T_326 = _T_317[7]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299356.4]
  assign _T_327 = _T_317[8]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299357.4]
  assign _T_328 = _T_317[9]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299358.4]
  assign _T_329 = _T_317[10]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299359.4]
  assign _T_330 = _T_317[11]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299360.4]
  assign _T_331 = _T_317[12]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299361.4]
  assign _T_332 = _T_317[13]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299362.4]
  assign _T_333 = _T_317[14]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299363.4]
  assign _T_334 = _T_317[15]; // @[UserYanker.scala 59:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299364.4]
  assign _T_335 = auto_out_r_valid & auto_in_r_ready; // @[UserYanker.scala 61:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299365.4]
  assign _T_336 = _T_335 & _T_319; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299366.4]
  assign _T_338 = auto_in_ar_valid & auto_out_ar_ready; // @[UserYanker.scala 62:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299369.4]
  assign _T_341 = _T_335 & _T_320; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299374.4]
  assign _T_346 = _T_335 & _T_321; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299382.4]
  assign _T_351 = _T_335 & _T_322; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299390.4]
  assign _T_356 = _T_335 & _T_323; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299398.4]
  assign _T_361 = _T_335 & _T_324; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299406.4]
  assign _T_366 = _T_335 & _T_325; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299414.4]
  assign _T_371 = _T_335 & _T_326; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299422.4]
  assign _T_376 = _T_335 & _T_327; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299430.4]
  assign _T_381 = _T_335 & _T_328; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299438.4]
  assign _T_386 = _T_335 & _T_329; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299446.4]
  assign _T_391 = _T_335 & _T_330; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299454.4]
  assign _T_396 = _T_335 & _T_331; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299462.4]
  assign _T_401 = _T_335 & _T_332; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299470.4]
  assign _T_406 = _T_335 & _T_333; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299478.4]
  assign _T_411 = _T_335 & _T_334; // @[UserYanker.scala 61:53:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299486.4]
  assign _T_418_0 = Queue_16_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299495.4]
  assign _T_418_1 = Queue_17_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299496.4]
  assign _GEN_49 = 4'h1 == auto_in_aw_bits_id ? _T_418_1 : _T_418_0; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_2 = Queue_18_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299497.4]
  assign _GEN_50 = 4'h2 == auto_in_aw_bits_id ? _T_418_2 : _GEN_49; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_3 = Queue_19_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299498.4]
  assign _GEN_51 = 4'h3 == auto_in_aw_bits_id ? _T_418_3 : _GEN_50; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_4 = Queue_20_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299499.4]
  assign _GEN_52 = 4'h4 == auto_in_aw_bits_id ? _T_418_4 : _GEN_51; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_5 = Queue_21_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299500.4]
  assign _GEN_53 = 4'h5 == auto_in_aw_bits_id ? _T_418_5 : _GEN_52; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_6 = Queue_22_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299501.4]
  assign _GEN_54 = 4'h6 == auto_in_aw_bits_id ? _T_418_6 : _GEN_53; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_7 = Queue_23_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299502.4]
  assign _GEN_55 = 4'h7 == auto_in_aw_bits_id ? _T_418_7 : _GEN_54; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_8 = Queue_24_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299503.4]
  assign _GEN_56 = 4'h8 == auto_in_aw_bits_id ? _T_418_8 : _GEN_55; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_9 = Queue_25_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299504.4]
  assign _GEN_57 = 4'h9 == auto_in_aw_bits_id ? _T_418_9 : _GEN_56; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_10 = Queue_26_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299505.4]
  assign _GEN_58 = 4'ha == auto_in_aw_bits_id ? _T_418_10 : _GEN_57; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_11 = Queue_27_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299506.4]
  assign _GEN_59 = 4'hb == auto_in_aw_bits_id ? _T_418_11 : _GEN_58; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_12 = Queue_28_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299507.4]
  assign _GEN_60 = 4'hc == auto_in_aw_bits_id ? _T_418_12 : _GEN_59; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_13 = Queue_29_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299508.4]
  assign _GEN_61 = 4'hd == auto_in_aw_bits_id ? _T_418_13 : _GEN_60; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_14 = Queue_30_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299509.4]
  assign _GEN_62 = 4'he == auto_in_aw_bits_id ? _T_418_14 : _GEN_61; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_418_15 = Queue_31_io_enq_ready; // @[UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299493.4 UserYanker.scala 67:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299510.4]
  assign _GEN_63 = 4'hf == auto_in_aw_bits_id ? _T_418_15 : _GEN_62; // @[UserYanker.scala 68:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299511.4]
  assign _T_486 = auto_out_b_valid == 1'h0; // @[UserYanker.scala 75:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299552.4]
  assign _T_443_0 = Queue_16_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299518.4]
  assign _T_443_1 = Queue_17_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299519.4]
  assign _GEN_65 = 4'h1 == auto_out_b_bits_id ? _T_443_1 : _T_443_0; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_2 = Queue_18_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299520.4]
  assign _GEN_66 = 4'h2 == auto_out_b_bits_id ? _T_443_2 : _GEN_65; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_3 = Queue_19_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299521.4]
  assign _GEN_67 = 4'h3 == auto_out_b_bits_id ? _T_443_3 : _GEN_66; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_4 = Queue_20_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299522.4]
  assign _GEN_68 = 4'h4 == auto_out_b_bits_id ? _T_443_4 : _GEN_67; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_5 = Queue_21_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299523.4]
  assign _GEN_69 = 4'h5 == auto_out_b_bits_id ? _T_443_5 : _GEN_68; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_6 = Queue_22_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299524.4]
  assign _GEN_70 = 4'h6 == auto_out_b_bits_id ? _T_443_6 : _GEN_69; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_7 = Queue_23_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299525.4]
  assign _GEN_71 = 4'h7 == auto_out_b_bits_id ? _T_443_7 : _GEN_70; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_8 = Queue_24_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299526.4]
  assign _GEN_72 = 4'h8 == auto_out_b_bits_id ? _T_443_8 : _GEN_71; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_9 = Queue_25_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299527.4]
  assign _GEN_73 = 4'h9 == auto_out_b_bits_id ? _T_443_9 : _GEN_72; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_10 = Queue_26_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299528.4]
  assign _GEN_74 = 4'ha == auto_out_b_bits_id ? _T_443_10 : _GEN_73; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_11 = Queue_27_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299529.4]
  assign _GEN_75 = 4'hb == auto_out_b_bits_id ? _T_443_11 : _GEN_74; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_12 = Queue_28_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299530.4]
  assign _GEN_76 = 4'hc == auto_out_b_bits_id ? _T_443_12 : _GEN_75; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_13 = Queue_29_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299531.4]
  assign _GEN_77 = 4'hd == auto_out_b_bits_id ? _T_443_13 : _GEN_76; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_14 = Queue_30_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299532.4]
  assign _GEN_78 = 4'he == auto_out_b_bits_id ? _T_443_14 : _GEN_77; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_443_15 = Queue_31_io_deq_valid; // @[UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299516.4 UserYanker.scala 73:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299533.4]
  assign _GEN_79 = 4'hf == auto_out_b_bits_id ? _T_443_15 : _GEN_78; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_487 = _T_486 | _GEN_79; // @[UserYanker.scala 75:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299553.4]
  assign _T_489 = _T_487 | reset; // @[UserYanker.scala 75:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299555.4]
  assign _T_490 = _T_489 == 1'h0; // @[UserYanker.scala 75:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299556.4]
  assign _T_466_0 = Queue_16_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299536.4]
  assign _T_466_1 = Queue_17_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299537.4]
  assign _GEN_81 = 4'h1 == auto_out_b_bits_id ? _T_466_1 : _T_466_0; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_2 = Queue_18_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299538.4]
  assign _GEN_82 = 4'h2 == auto_out_b_bits_id ? _T_466_2 : _GEN_81; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_3 = Queue_19_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299539.4]
  assign _GEN_83 = 4'h3 == auto_out_b_bits_id ? _T_466_3 : _GEN_82; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_4 = Queue_20_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299540.4]
  assign _GEN_84 = 4'h4 == auto_out_b_bits_id ? _T_466_4 : _GEN_83; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_5 = Queue_21_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299541.4]
  assign _GEN_85 = 4'h5 == auto_out_b_bits_id ? _T_466_5 : _GEN_84; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_6 = Queue_22_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299542.4]
  assign _GEN_86 = 4'h6 == auto_out_b_bits_id ? _T_466_6 : _GEN_85; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_7 = Queue_23_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299543.4]
  assign _GEN_87 = 4'h7 == auto_out_b_bits_id ? _T_466_7 : _GEN_86; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_8 = Queue_24_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299544.4]
  assign _GEN_88 = 4'h8 == auto_out_b_bits_id ? _T_466_8 : _GEN_87; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_9 = Queue_25_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299545.4]
  assign _GEN_89 = 4'h9 == auto_out_b_bits_id ? _T_466_9 : _GEN_88; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_10 = Queue_26_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299546.4]
  assign _GEN_90 = 4'ha == auto_out_b_bits_id ? _T_466_10 : _GEN_89; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_11 = Queue_27_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299547.4]
  assign _GEN_91 = 4'hb == auto_out_b_bits_id ? _T_466_11 : _GEN_90; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_12 = Queue_28_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299548.4]
  assign _GEN_92 = 4'hc == auto_out_b_bits_id ? _T_466_12 : _GEN_91; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_13 = Queue_29_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299549.4]
  assign _GEN_93 = 4'hd == auto_out_b_bits_id ? _T_466_13 : _GEN_92; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_14 = Queue_30_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299550.4]
  assign _GEN_94 = 4'he == auto_out_b_bits_id ? _T_466_14 : _GEN_93; // @[UserYanker.scala 77:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299562.4]
  assign _T_466_15 = Queue_31_io_deq_bits; // @[UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299534.4 UserYanker.scala 74:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299551.4]
  assign _T_492 = 16'h1 << auto_in_aw_bits_id; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299564.4]
  assign _T_494 = _T_492[0]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299566.4]
  assign _T_495 = _T_492[1]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299567.4]
  assign _T_496 = _T_492[2]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299568.4]
  assign _T_497 = _T_492[3]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299569.4]
  assign _T_498 = _T_492[4]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299570.4]
  assign _T_499 = _T_492[5]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299571.4]
  assign _T_500 = _T_492[6]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299572.4]
  assign _T_501 = _T_492[7]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299573.4]
  assign _T_502 = _T_492[8]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299574.4]
  assign _T_503 = _T_492[9]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299575.4]
  assign _T_504 = _T_492[10]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299576.4]
  assign _T_505 = _T_492[11]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299577.4]
  assign _T_506 = _T_492[12]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299578.4]
  assign _T_507 = _T_492[13]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299579.4]
  assign _T_508 = _T_492[14]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299580.4]
  assign _T_509 = _T_492[15]; // @[UserYanker.scala 79:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299581.4]
  assign _T_511 = 16'h1 << auto_out_b_bits_id; // @[OneHot.scala 52:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299583.4]
  assign _T_513 = _T_511[0]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299585.4]
  assign _T_514 = _T_511[1]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299586.4]
  assign _T_515 = _T_511[2]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299587.4]
  assign _T_516 = _T_511[3]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299588.4]
  assign _T_517 = _T_511[4]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299589.4]
  assign _T_518 = _T_511[5]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299590.4]
  assign _T_519 = _T_511[6]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299591.4]
  assign _T_520 = _T_511[7]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299592.4]
  assign _T_521 = _T_511[8]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299593.4]
  assign _T_522 = _T_511[9]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299594.4]
  assign _T_523 = _T_511[10]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299595.4]
  assign _T_524 = _T_511[11]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299596.4]
  assign _T_525 = _T_511[12]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299597.4]
  assign _T_526 = _T_511[13]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299598.4]
  assign _T_527 = _T_511[14]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299599.4]
  assign _T_528 = _T_511[15]; // @[UserYanker.scala 80:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299600.4]
  assign _T_529 = auto_out_b_valid & auto_in_b_ready; // @[UserYanker.scala 82:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299601.4]
  assign _T_531 = auto_in_aw_valid & auto_out_aw_ready; // @[UserYanker.scala 83:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299604.4]
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_63; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_b_bits_user = 4'hf == auto_out_b_bits_id ? _T_466_15 : _GEN_94; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_15; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_r_bits_user = 4'hf == auto_out_r_bits_id ? _T_272_15 : _GEN_46; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299128.4]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_63; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_15; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299127.4]
  assign Queue_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299131.4]
  assign Queue_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299132.4]
  assign Queue_io_enq_valid = _T_338 & _T_300; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299371.4]
  assign Queue_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299372.4]
  assign Queue_io_deq_ready = _T_336 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299368.4]
  assign Queue_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299135.4]
  assign Queue_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299136.4]
  assign Queue_1_io_enq_valid = _T_338 & _T_301; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299379.4]
  assign Queue_1_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299380.4]
  assign Queue_1_io_deq_ready = _T_341 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299376.4]
  assign Queue_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299139.4]
  assign Queue_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299140.4]
  assign Queue_2_io_enq_valid = _T_338 & _T_302; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299387.4]
  assign Queue_2_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299388.4]
  assign Queue_2_io_deq_ready = _T_346 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299384.4]
  assign Queue_3_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299143.4]
  assign Queue_3_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299144.4]
  assign Queue_3_io_enq_valid = _T_338 & _T_303; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299395.4]
  assign Queue_3_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299396.4]
  assign Queue_3_io_deq_ready = _T_351 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299392.4]
  assign Queue_4_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299147.4]
  assign Queue_4_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299148.4]
  assign Queue_4_io_enq_valid = _T_338 & _T_304; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299403.4]
  assign Queue_4_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299404.4]
  assign Queue_4_io_deq_ready = _T_356 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299400.4]
  assign Queue_5_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299151.4]
  assign Queue_5_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299152.4]
  assign Queue_5_io_enq_valid = _T_338 & _T_305; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299411.4]
  assign Queue_5_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299412.4]
  assign Queue_5_io_deq_ready = _T_361 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299408.4]
  assign Queue_6_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299155.4]
  assign Queue_6_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299156.4]
  assign Queue_6_io_enq_valid = _T_338 & _T_306; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299419.4]
  assign Queue_6_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299420.4]
  assign Queue_6_io_deq_ready = _T_366 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299416.4]
  assign Queue_7_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299159.4]
  assign Queue_7_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299160.4]
  assign Queue_7_io_enq_valid = _T_338 & _T_307; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299427.4]
  assign Queue_7_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299428.4]
  assign Queue_7_io_deq_ready = _T_371 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299424.4]
  assign Queue_8_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299163.4]
  assign Queue_8_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299164.4]
  assign Queue_8_io_enq_valid = _T_338 & _T_308; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299435.4]
  assign Queue_8_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299436.4]
  assign Queue_8_io_deq_ready = _T_376 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299432.4]
  assign Queue_9_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299167.4]
  assign Queue_9_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299168.4]
  assign Queue_9_io_enq_valid = _T_338 & _T_309; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299443.4]
  assign Queue_9_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299444.4]
  assign Queue_9_io_deq_ready = _T_381 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299440.4]
  assign Queue_10_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299171.4]
  assign Queue_10_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299172.4]
  assign Queue_10_io_enq_valid = _T_338 & _T_310; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299451.4]
  assign Queue_10_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299452.4]
  assign Queue_10_io_deq_ready = _T_386 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299448.4]
  assign Queue_11_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299175.4]
  assign Queue_11_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299176.4]
  assign Queue_11_io_enq_valid = _T_338 & _T_311; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299459.4]
  assign Queue_11_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299460.4]
  assign Queue_11_io_deq_ready = _T_391 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299456.4]
  assign Queue_12_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299179.4]
  assign Queue_12_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299180.4]
  assign Queue_12_io_enq_valid = _T_338 & _T_312; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299467.4]
  assign Queue_12_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299468.4]
  assign Queue_12_io_deq_ready = _T_396 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299464.4]
  assign Queue_13_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299183.4]
  assign Queue_13_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299184.4]
  assign Queue_13_io_enq_valid = _T_338 & _T_313; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299475.4]
  assign Queue_13_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299476.4]
  assign Queue_13_io_deq_ready = _T_401 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299472.4]
  assign Queue_14_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299187.4]
  assign Queue_14_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299188.4]
  assign Queue_14_io_enq_valid = _T_338 & _T_314; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299483.4]
  assign Queue_14_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299484.4]
  assign Queue_14_io_deq_ready = _T_406 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299480.4]
  assign Queue_15_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299191.4]
  assign Queue_15_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299192.4]
  assign Queue_15_io_enq_valid = _T_338 & _T_315; // @[UserYanker.scala 62:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299491.4]
  assign Queue_15_io_enq_bits = auto_in_ar_bits_user; // @[UserYanker.scala 63:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299492.4]
  assign Queue_15_io_deq_ready = _T_411 & auto_out_r_bits_last; // @[UserYanker.scala 61:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299488.4]
  assign Queue_16_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299195.4]
  assign Queue_16_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299196.4]
  assign Queue_16_io_enq_valid = _T_531 & _T_494; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299606.4]
  assign Queue_16_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299607.4]
  assign Queue_16_io_deq_ready = _T_529 & _T_513; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299603.4]
  assign Queue_17_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299199.4]
  assign Queue_17_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299200.4]
  assign Queue_17_io_enq_valid = _T_531 & _T_495; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299613.4]
  assign Queue_17_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299614.4]
  assign Queue_17_io_deq_ready = _T_529 & _T_514; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299610.4]
  assign Queue_18_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299203.4]
  assign Queue_18_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299204.4]
  assign Queue_18_io_enq_valid = _T_531 & _T_496; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299620.4]
  assign Queue_18_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299621.4]
  assign Queue_18_io_deq_ready = _T_529 & _T_515; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299617.4]
  assign Queue_19_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299207.4]
  assign Queue_19_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299208.4]
  assign Queue_19_io_enq_valid = _T_531 & _T_497; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299627.4]
  assign Queue_19_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299628.4]
  assign Queue_19_io_deq_ready = _T_529 & _T_516; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299624.4]
  assign Queue_20_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299211.4]
  assign Queue_20_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299212.4]
  assign Queue_20_io_enq_valid = _T_531 & _T_498; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299634.4]
  assign Queue_20_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299635.4]
  assign Queue_20_io_deq_ready = _T_529 & _T_517; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299631.4]
  assign Queue_21_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299215.4]
  assign Queue_21_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299216.4]
  assign Queue_21_io_enq_valid = _T_531 & _T_499; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299641.4]
  assign Queue_21_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299642.4]
  assign Queue_21_io_deq_ready = _T_529 & _T_518; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299638.4]
  assign Queue_22_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299219.4]
  assign Queue_22_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299220.4]
  assign Queue_22_io_enq_valid = _T_531 & _T_500; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299648.4]
  assign Queue_22_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299649.4]
  assign Queue_22_io_deq_ready = _T_529 & _T_519; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299645.4]
  assign Queue_23_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299223.4]
  assign Queue_23_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299224.4]
  assign Queue_23_io_enq_valid = _T_531 & _T_501; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299655.4]
  assign Queue_23_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299656.4]
  assign Queue_23_io_deq_ready = _T_529 & _T_520; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299652.4]
  assign Queue_24_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299227.4]
  assign Queue_24_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299228.4]
  assign Queue_24_io_enq_valid = _T_531 & _T_502; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299662.4]
  assign Queue_24_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299663.4]
  assign Queue_24_io_deq_ready = _T_529 & _T_521; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299659.4]
  assign Queue_25_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299231.4]
  assign Queue_25_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299232.4]
  assign Queue_25_io_enq_valid = _T_531 & _T_503; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299669.4]
  assign Queue_25_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299670.4]
  assign Queue_25_io_deq_ready = _T_529 & _T_522; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299666.4]
  assign Queue_26_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299235.4]
  assign Queue_26_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299236.4]
  assign Queue_26_io_enq_valid = _T_531 & _T_504; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299676.4]
  assign Queue_26_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299677.4]
  assign Queue_26_io_deq_ready = _T_529 & _T_523; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299673.4]
  assign Queue_27_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299239.4]
  assign Queue_27_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299240.4]
  assign Queue_27_io_enq_valid = _T_531 & _T_505; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299683.4]
  assign Queue_27_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299684.4]
  assign Queue_27_io_deq_ready = _T_529 & _T_524; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299680.4]
  assign Queue_28_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299243.4]
  assign Queue_28_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299244.4]
  assign Queue_28_io_enq_valid = _T_531 & _T_506; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299690.4]
  assign Queue_28_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299691.4]
  assign Queue_28_io_deq_ready = _T_529 & _T_525; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299687.4]
  assign Queue_29_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299247.4]
  assign Queue_29_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299248.4]
  assign Queue_29_io_enq_valid = _T_531 & _T_507; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299697.4]
  assign Queue_29_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299698.4]
  assign Queue_29_io_deq_ready = _T_529 & _T_526; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299694.4]
  assign Queue_30_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299251.4]
  assign Queue_30_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299252.4]
  assign Queue_30_io_enq_valid = _T_531 & _T_508; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299704.4]
  assign Queue_30_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299705.4]
  assign Queue_30_io_deq_ready = _T_529 & _T_527; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299701.4]
  assign Queue_31_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299255.4]
  assign Queue_31_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299256.4]
  assign Queue_31_io_enq_valid = _T_531 & _T_509; // @[UserYanker.scala 83:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299711.4]
  assign Queue_31_io_enq_bits = auto_in_aw_bits_user; // @[UserYanker.scala 84:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299712.4]
  assign Queue_31_io_deq_ready = _T_529 & _T_528; // @[UserYanker.scala 82:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299708.4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_296) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:54 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"); // @[UserYanker.scala 54:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299322.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_296) begin
          $fatal; // @[UserYanker.scala 54:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299323.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_490) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:75 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"); // @[UserYanker.scala 75:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299558.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_490) begin
          $fatal; // @[UserYanker.scala 75:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@299559.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AsyncResetSynchronizerShiftReg_w4_d3_i0( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300103.2]
  input        clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300104.4]
  input        reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300105.4]
  input  [3:0] io_d, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300106.4]
  output [3:0] io_q // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300106.4]
);
  wire  sync_0_clock; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300111.4]
  wire  sync_0_reset; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300111.4]
  wire [3:0] sync_0_io_d; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300111.4]
  wire [3:0] sync_0_io_q; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300111.4]
  wire  sync_0_io_en; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300111.4]
  wire  sync_1_clock; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300115.4]
  wire  sync_1_reset; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300115.4]
  wire [3:0] sync_1_io_d; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300115.4]
  wire [3:0] sync_1_io_q; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300115.4]
  wire  sync_1_io_en; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300115.4]
  wire  sync_2_clock; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300119.4]
  wire  sync_2_reset; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300119.4]
  wire [3:0] sync_2_io_d; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300119.4]
  wire [3:0] sync_2_io_q; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300119.4]
  wire  sync_2_io_en; // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300119.4]
  AsyncResetRegVec_w4_i0 sync_0 ( // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300111.4]
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  AsyncResetRegVec_w4_i0 sync_1 ( // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300115.4]
    .clock(sync_1_clock),
    .reset(sync_1_reset),
    .io_d(sync_1_io_d),
    .io_q(sync_1_io_q),
    .io_en(sync_1_io_en)
  );
  AsyncResetRegVec_w4_i0 sync_2 ( // @[ShiftReg.scala 60:12:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300119.4]
    .clock(sync_2_clock),
    .reset(sync_2_reset),
    .io_d(sync_2_io_d),
    .io_q(sync_2_io_q),
    .io_en(sync_2_io_en)
  );
  assign io_q = sync_0_io_q; // @[ShiftReg.scala 70:8:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300129.4]
  assign sync_0_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300113.4]
  assign sync_0_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300114.4]
  assign sync_0_io_d = sync_1_io_q; // @[ShiftReg.scala 67:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300125.4]
  assign sync_0_io_en = 1'h1; // @[ShiftReg.scala 68:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300126.4]
  assign sync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300117.4]
  assign sync_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300118.4]
  assign sync_1_io_d = sync_2_io_q; // @[ShiftReg.scala 67:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300127.4]
  assign sync_1_io_en = 1'h1; // @[ShiftReg.scala 68:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300128.4]
  assign sync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300121.4]
  assign sync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300122.4]
  assign sync_2_io_d = io_d; // @[ShiftReg.scala 63:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300123.4]
  assign sync_2_io_en = 1'h1; // @[ShiftReg.scala 64:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300124.4]
endmodule
module SynchronizerShiftReg_w61_d1( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300131.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300132.4]
  input  [60:0] io_d, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300134.4]
  output [60:0] io_q // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300134.4]
);
  reg [60:0] sync_0; // @[ShiftReg.scala 114:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300139.4]
  reg [63:0] _RAND_0;
  assign io_q = sync_0; // @[ShiftReg.scala 123:8:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300141.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  sync_0 = _RAND_0[60:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    sync_0 <= io_d;
  end
endmodule
module AsyncQueueSink_3( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300673.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300674.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300675.4]
  input         io_deq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output        io_deq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [3:0]  io_deq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [31:0] io_deq_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [7:0]  io_deq_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [2:0]  io_deq_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [1:0]  io_deq_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output        io_deq_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [3:0]  io_deq_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [2:0]  io_deq_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [3:0]  io_deq_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [31:0] io_async_mem_0_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [7:0]  io_async_mem_0_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_0_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [1:0]  io_async_mem_0_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_mem_0_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_0_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_0_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_0_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [31:0] io_async_mem_1_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [7:0]  io_async_mem_1_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_1_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [1:0]  io_async_mem_1_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_mem_1_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_1_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_1_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_1_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [31:0] io_async_mem_2_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [7:0]  io_async_mem_2_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_2_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [1:0]  io_async_mem_2_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_mem_2_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_2_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_2_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_2_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [31:0] io_async_mem_3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [7:0]  io_async_mem_3_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_3_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [1:0]  io_async_mem_3_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_mem_3_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_3_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_3_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_3_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [31:0] io_async_mem_4_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [7:0]  io_async_mem_4_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_4_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [1:0]  io_async_mem_4_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_mem_4_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_4_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_4_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_4_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [31:0] io_async_mem_5_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [7:0]  io_async_mem_5_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_5_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [1:0]  io_async_mem_5_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_mem_5_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_5_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_5_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_5_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [31:0] io_async_mem_6_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [7:0]  io_async_mem_6_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_6_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [1:0]  io_async_mem_6_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_mem_6_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_6_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_6_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_6_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [31:0] io_async_mem_7_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [7:0]  io_async_mem_7_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_7_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [1:0]  io_async_mem_7_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_mem_7_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_7_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [2:0]  io_async_mem_7_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_mem_7_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output [3:0]  io_async_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input  [3:0]  io_async_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output        io_async_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  input         io_async_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
  output        io_async_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300676.4]
);
  wire  ridx_bin_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300683.4]
  wire  ridx_bin_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300683.4]
  wire [3:0] ridx_bin_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300683.4]
  wire [3:0] ridx_bin_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300683.4]
  wire  ridx_bin_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300683.4]
  wire  widx_gray_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300695.4]
  wire  widx_gray_reset; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300695.4]
  wire [3:0] widx_gray_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300695.4]
  wire [3:0] widx_gray_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300695.4]
  wire  deq_bits_reg_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300710.4]
  wire [60:0] deq_bits_reg_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300710.4]
  wire [60:0] deq_bits_reg_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300710.4]
  wire  valid_reg_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300755.4]
  wire  valid_reg_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300755.4]
  wire  valid_reg_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300755.4]
  wire  valid_reg_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300755.4]
  wire  valid_reg_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300755.4]
  wire  ridx_gray_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300764.4]
  wire  ridx_gray_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300764.4]
  wire [3:0] ridx_gray_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300764.4]
  wire [3:0] ridx_gray_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300764.4]
  wire  ridx_gray_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300764.4]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300771.4]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300771.4]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300771.4]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300771.4]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300774.4]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300774.4]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300774.4]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300774.4]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300777.4]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300777.4]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300777.4]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300777.4]
  wire  AsyncResetRegVec_w1_i0_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300806.4]
  wire  AsyncResetRegVec_w1_i0_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300806.4]
  wire  AsyncResetRegVec_w1_i0_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300806.4]
  wire  AsyncResetRegVec_w1_i0_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300806.4]
  wire  AsyncResetRegVec_w1_i0_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300806.4]
  wire  _T_86; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300680.4]
  wire  source_ready; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300678.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300679.4 AsyncQueue.scala 164:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300792.4]
  wire  _T_87; // @[AsyncQueue.scala 130:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300681.4]
  wire [3:0] _GEN_72; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300689.4]
  wire [3:0] _T_91; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300690.4]
  wire [3:0] _T_92; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300691.4]
  wire [2:0] _T_93; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300693.4]
  wire [3:0] _GEN_73; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300694.4]
  wire [3:0] ridx; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300694.4]
  wire [3:0] widx; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300700.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300702.4]
  wire  _T_95; // @[AsyncQueue.scala 132:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300703.4]
  wire  valid; // @[AsyncQueue.scala 132:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300704.4]
  wire [2:0] _T_96; // @[AsyncQueue.scala 138:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300705.4]
  wire  _T_97; // @[AsyncQueue.scala 138:62:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300706.4]
  wire [2:0] _GEN_74; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300707.4]
  wire [2:0] _T_98; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300707.4]
  wire [2:0] index; // @[AsyncQueue.scala 138:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300708.4]
  wire [3:0] _GEN_9; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [31:0] _GEN_10; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [7:0] _GEN_11; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_12; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [1:0] _GEN_13; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire  _GEN_14; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_15; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_16; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_17; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_18; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [31:0] _GEN_19; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [7:0] _GEN_20; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_21; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [1:0] _GEN_22; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire  _GEN_23; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_24; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_25; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_26; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_27; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [31:0] _GEN_28; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [7:0] _GEN_29; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_30; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [1:0] _GEN_31; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire  _GEN_32; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_33; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_34; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_35; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_36; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [31:0] _GEN_37; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [7:0] _GEN_38; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_39; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [1:0] _GEN_40; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire  _GEN_41; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_42; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_43; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_44; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_45; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [31:0] _GEN_46; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [7:0] _GEN_47; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_48; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [1:0] _GEN_49; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire  _GEN_50; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_51; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_52; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_53; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_54; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [31:0] _GEN_55; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [7:0] _GEN_56; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_57; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [1:0] _GEN_58; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire  _GEN_59; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_60; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_61; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_62; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_63; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [31:0] _GEN_64; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [7:0] _GEN_65; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_66; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [1:0] _GEN_67; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire  _GEN_68; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_69; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] _GEN_70; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] _GEN_71; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] deq_bits_nxt_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [31:0] deq_bits_nxt_addr; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [7:0] deq_bits_nxt_len; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] deq_bits_nxt_size; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [1:0] deq_bits_nxt_burst; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire  deq_bits_nxt_lock; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] deq_bits_nxt_cache; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [2:0] deq_bits_nxt_prot; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [3:0] deq_bits_nxt_qos; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  wire [6:0] _T_100; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300714.4]
  wire [4:0] _T_101; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300715.4]
  wire [11:0] _T_102; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300716.4]
  wire [4:0] _T_103; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300717.4]
  wire [35:0] _T_104; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300718.4]
  wire [43:0] _T_105; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300719.4]
  wire [48:0] _T_106; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300720.4]
  wire [60:0] _T_111; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300725.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300727.4]
  wire  valid_reg_1; // @[AsyncQueue.scala 147:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300761.4]
  wire  _T_123; // @[AsyncQueue.scala 157:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300781.4]
  AsyncResetRegVec_w4_i0 ridx_bin ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300683.4]
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_gray ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300695.4]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  SynchronizerShiftReg_w61_d1 deq_bits_reg ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300710.4]
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q)
  );
  AsyncResetRegVec_w1_i0 valid_reg ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300755.4]
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_w4_i0 ridx_gray ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300764.4]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300771.4]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300774.4]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300777.4]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300806.4]
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q),
    .io_en(AsyncResetRegVec_w1_i0_io_en)
  );
  assign _T_86 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300680.4]
  assign source_ready = AsyncValidSync_2_io_out; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300678.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300679.4 AsyncQueue.scala 164:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300792.4]
  assign _T_87 = source_ready == 1'h0; // @[AsyncQueue.scala 130:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300681.4]
  assign _GEN_72 = {{3'd0}, _T_86}; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300689.4]
  assign _T_91 = ridx_bin_io_q + _GEN_72; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300690.4]
  assign _T_92 = _T_87 ? 4'h0 : _T_91; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300691.4]
  assign _T_93 = _T_92[3:1]; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300693.4]
  assign _GEN_73 = {{1'd0}, _T_93}; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300694.4]
  assign ridx = _T_92 ^ _GEN_73; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300694.4]
  assign widx = widx_gray_io_q; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300700.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300702.4]
  assign _T_95 = ridx != widx; // @[AsyncQueue.scala 132:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300703.4]
  assign valid = source_ready & _T_95; // @[AsyncQueue.scala 132:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300704.4]
  assign _T_96 = ridx[2:0]; // @[AsyncQueue.scala 138:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300705.4]
  assign _T_97 = ridx[3]; // @[AsyncQueue.scala 138:62:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300706.4]
  assign _GEN_74 = {{2'd0}, _T_97}; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300707.4]
  assign _T_98 = _GEN_74 << 2; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300707.4]
  assign index = _T_96 ^ _T_98; // @[AsyncQueue.scala 138:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300708.4]
  assign _GEN_9 = 3'h1 == index ? io_async_mem_1_id : io_async_mem_0_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_10 = 3'h1 == index ? io_async_mem_1_addr : io_async_mem_0_addr; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_11 = 3'h1 == index ? io_async_mem_1_len : io_async_mem_0_len; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_12 = 3'h1 == index ? io_async_mem_1_size : io_async_mem_0_size; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_13 = 3'h1 == index ? io_async_mem_1_burst : io_async_mem_0_burst; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_14 = 3'h1 == index ? io_async_mem_1_lock : io_async_mem_0_lock; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_15 = 3'h1 == index ? io_async_mem_1_cache : io_async_mem_0_cache; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_16 = 3'h1 == index ? io_async_mem_1_prot : io_async_mem_0_prot; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_17 = 3'h1 == index ? io_async_mem_1_qos : io_async_mem_0_qos; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_18 = 3'h2 == index ? io_async_mem_2_id : _GEN_9; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_19 = 3'h2 == index ? io_async_mem_2_addr : _GEN_10; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_20 = 3'h2 == index ? io_async_mem_2_len : _GEN_11; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_21 = 3'h2 == index ? io_async_mem_2_size : _GEN_12; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_22 = 3'h2 == index ? io_async_mem_2_burst : _GEN_13; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_23 = 3'h2 == index ? io_async_mem_2_lock : _GEN_14; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_24 = 3'h2 == index ? io_async_mem_2_cache : _GEN_15; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_25 = 3'h2 == index ? io_async_mem_2_prot : _GEN_16; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_26 = 3'h2 == index ? io_async_mem_2_qos : _GEN_17; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_27 = 3'h3 == index ? io_async_mem_3_id : _GEN_18; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_28 = 3'h3 == index ? io_async_mem_3_addr : _GEN_19; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_29 = 3'h3 == index ? io_async_mem_3_len : _GEN_20; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_30 = 3'h3 == index ? io_async_mem_3_size : _GEN_21; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_31 = 3'h3 == index ? io_async_mem_3_burst : _GEN_22; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_32 = 3'h3 == index ? io_async_mem_3_lock : _GEN_23; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_33 = 3'h3 == index ? io_async_mem_3_cache : _GEN_24; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_34 = 3'h3 == index ? io_async_mem_3_prot : _GEN_25; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_35 = 3'h3 == index ? io_async_mem_3_qos : _GEN_26; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_36 = 3'h4 == index ? io_async_mem_4_id : _GEN_27; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_37 = 3'h4 == index ? io_async_mem_4_addr : _GEN_28; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_38 = 3'h4 == index ? io_async_mem_4_len : _GEN_29; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_39 = 3'h4 == index ? io_async_mem_4_size : _GEN_30; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_40 = 3'h4 == index ? io_async_mem_4_burst : _GEN_31; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_41 = 3'h4 == index ? io_async_mem_4_lock : _GEN_32; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_42 = 3'h4 == index ? io_async_mem_4_cache : _GEN_33; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_43 = 3'h4 == index ? io_async_mem_4_prot : _GEN_34; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_44 = 3'h4 == index ? io_async_mem_4_qos : _GEN_35; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_45 = 3'h5 == index ? io_async_mem_5_id : _GEN_36; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_46 = 3'h5 == index ? io_async_mem_5_addr : _GEN_37; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_47 = 3'h5 == index ? io_async_mem_5_len : _GEN_38; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_48 = 3'h5 == index ? io_async_mem_5_size : _GEN_39; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_49 = 3'h5 == index ? io_async_mem_5_burst : _GEN_40; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_50 = 3'h5 == index ? io_async_mem_5_lock : _GEN_41; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_51 = 3'h5 == index ? io_async_mem_5_cache : _GEN_42; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_52 = 3'h5 == index ? io_async_mem_5_prot : _GEN_43; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_53 = 3'h5 == index ? io_async_mem_5_qos : _GEN_44; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_54 = 3'h6 == index ? io_async_mem_6_id : _GEN_45; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_55 = 3'h6 == index ? io_async_mem_6_addr : _GEN_46; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_56 = 3'h6 == index ? io_async_mem_6_len : _GEN_47; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_57 = 3'h6 == index ? io_async_mem_6_size : _GEN_48; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_58 = 3'h6 == index ? io_async_mem_6_burst : _GEN_49; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_59 = 3'h6 == index ? io_async_mem_6_lock : _GEN_50; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_60 = 3'h6 == index ? io_async_mem_6_cache : _GEN_51; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_61 = 3'h6 == index ? io_async_mem_6_prot : _GEN_52; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_62 = 3'h6 == index ? io_async_mem_6_qos : _GEN_53; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_63 = 3'h7 == index ? io_async_mem_7_id : _GEN_54; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_64 = 3'h7 == index ? io_async_mem_7_addr : _GEN_55; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_65 = 3'h7 == index ? io_async_mem_7_len : _GEN_56; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_66 = 3'h7 == index ? io_async_mem_7_size : _GEN_57; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_67 = 3'h7 == index ? io_async_mem_7_burst : _GEN_58; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_68 = 3'h7 == index ? io_async_mem_7_lock : _GEN_59; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_69 = 3'h7 == index ? io_async_mem_7_cache : _GEN_60; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_70 = 3'h7 == index ? io_async_mem_7_prot : _GEN_61; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _GEN_71 = 3'h7 == index ? io_async_mem_7_qos : _GEN_62; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_id = valid ? _GEN_63 : io_deq_bits_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_addr = valid ? _GEN_64 : io_deq_bits_addr; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_len = valid ? _GEN_65 : io_deq_bits_len; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_size = valid ? _GEN_66 : io_deq_bits_size; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_burst = valid ? _GEN_67 : io_deq_bits_burst; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_lock = valid ? _GEN_68 : io_deq_bits_lock; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_cache = valid ? _GEN_69 : io_deq_bits_cache; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_prot = valid ? _GEN_70 : io_deq_bits_prot; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign deq_bits_nxt_qos = valid ? _GEN_71 : io_deq_bits_qos; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300709.4]
  assign _T_100 = {deq_bits_nxt_prot,deq_bits_nxt_qos}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300714.4]
  assign _T_101 = {deq_bits_nxt_lock,deq_bits_nxt_cache}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300715.4]
  assign _T_102 = {_T_101,_T_100}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300716.4]
  assign _T_103 = {deq_bits_nxt_size,deq_bits_nxt_burst}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300717.4]
  assign _T_104 = {deq_bits_nxt_id,deq_bits_nxt_addr}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300718.4]
  assign _T_105 = {_T_104,deq_bits_nxt_len}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300719.4]
  assign _T_106 = {_T_105,_T_103}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300720.4]
  assign _T_111 = deq_bits_reg_io_q; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300725.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300727.4]
  assign valid_reg_1 = valid_reg_io_q; // @[AsyncQueue.scala 147:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300761.4]
  assign _T_123 = io_async_safe_source_reset_n == 1'h0; // @[AsyncQueue.scala 157:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300781.4]
  assign io_deq_valid = valid_reg_1 & source_ready; // @[AsyncQueue.scala 148:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300763.4]
  assign io_deq_bits_id = _T_111[60:57]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300754.4]
  assign io_deq_bits_addr = _T_111[56:25]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300753.4]
  assign io_deq_bits_len = _T_111[24:17]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300752.4]
  assign io_deq_bits_size = _T_111[16:14]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300751.4]
  assign io_deq_bits_burst = _T_111[13:12]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300750.4]
  assign io_deq_bits_lock = _T_111[11]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300749.4]
  assign io_deq_bits_cache = _T_111[10:7]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300748.4]
  assign io_deq_bits_prot = _T_111[6:4]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300747.4]
  assign io_deq_bits_qos = _T_111[3:0]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300746.4]
  assign io_async_ridx = ridx_gray_io_q; // @[AsyncQueue.scala 151:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300770.4]
  assign io_async_safe_ridx_valid = AsyncValidSync_io_out; // @[AsyncQueue.scala 161:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300789.4]
  assign io_async_safe_sink_reset_n = reset == 1'h0; // @[AsyncQueue.scala 165:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300795.4]
  assign ridx_bin_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300685.4]
  assign ridx_bin_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300686.4]
  assign ridx_bin_io_d = _T_87 ? 4'h0 : _T_91; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300687.4]
  assign ridx_bin_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300688.4]
  assign widx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300697.4]
  assign widx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300698.4]
  assign widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300699.4]
  assign deq_bits_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300712.4]
  assign deq_bits_reg_io_d = {_T_106,_T_102}; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300722.4]
  assign valid_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300757.4]
  assign valid_reg_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300758.4]
  assign valid_reg_io_d = source_ready & _T_95; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300759.4]
  assign valid_reg_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300760.4]
  assign ridx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300766.4]
  assign ridx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300767.4]
  assign ridx_gray_io_d = _T_92 ^ _GEN_73; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300768.4]
  assign ridx_gray_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300769.4]
  assign AsyncValidSync_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300772.4]
  assign AsyncValidSync_reset = reset | _T_123; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300773.4 AsyncQueue.scala 157:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300783.4]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 160:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300788.4]
  assign AsyncValidSync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300775.4]
  assign AsyncValidSync_1_reset = reset | _T_123; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300776.4 AsyncQueue.scala 158:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300787.4]
  assign AsyncValidSync_1_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 162:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300790.4]
  assign AsyncValidSync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300778.4]
  assign AsyncValidSync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300779.4]
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 163:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300791.4]
  assign AsyncResetRegVec_w1_i0_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300808.4]
  assign AsyncResetRegVec_w1_i0_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300809.4]
  assign AsyncResetRegVec_w1_i0_io_d = io_async_widx == io_async_ridx; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300810.4]
  assign AsyncResetRegVec_w1_i0_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@300811.4]
endmodule
module SynchronizerShiftReg_w73_d1( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302327.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302328.4]
  input  [72:0] io_d, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302330.4]
  output [72:0] io_q // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302330.4]
);
  reg [72:0] sync_0; // @[ShiftReg.scala 114:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302335.4]
  reg [95:0] _RAND_0;
  assign io_q = sync_0; // @[ShiftReg.scala 123:8:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302337.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  sync_0 = _RAND_0[72:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    sync_0 <= io_d;
  end
endmodule
module AsyncQueueSink_5( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302869.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302870.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302871.4]
  input         io_deq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  output        io_deq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  output [63:0] io_deq_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  output [7:0]  io_deq_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  output        io_deq_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [63:0] io_async_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [7:0]  io_async_mem_0_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [63:0] io_async_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [7:0]  io_async_mem_1_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [63:0] io_async_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [7:0]  io_async_mem_2_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [63:0] io_async_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [7:0]  io_async_mem_3_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [63:0] io_async_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [7:0]  io_async_mem_4_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [63:0] io_async_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [7:0]  io_async_mem_5_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [63:0] io_async_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [7:0]  io_async_mem_6_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [63:0] io_async_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [7:0]  io_async_mem_7_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  output [3:0]  io_async_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input  [3:0]  io_async_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  output        io_async_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  input         io_async_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
  output        io_async_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302872.4]
);
  wire  ridx_bin_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302879.4]
  wire  ridx_bin_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302879.4]
  wire [3:0] ridx_bin_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302879.4]
  wire [3:0] ridx_bin_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302879.4]
  wire  ridx_bin_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302879.4]
  wire  widx_gray_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302891.4]
  wire  widx_gray_reset; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302891.4]
  wire [3:0] widx_gray_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302891.4]
  wire [3:0] widx_gray_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302891.4]
  wire  deq_bits_reg_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302906.4]
  wire [72:0] deq_bits_reg_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302906.4]
  wire [72:0] deq_bits_reg_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302906.4]
  wire  valid_reg_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302927.4]
  wire  valid_reg_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302927.4]
  wire  valid_reg_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302927.4]
  wire  valid_reg_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302927.4]
  wire  valid_reg_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302927.4]
  wire  ridx_gray_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302936.4]
  wire  ridx_gray_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302936.4]
  wire [3:0] ridx_gray_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302936.4]
  wire [3:0] ridx_gray_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302936.4]
  wire  ridx_gray_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302936.4]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302943.4]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302943.4]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302943.4]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302943.4]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302946.4]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302946.4]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302946.4]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302946.4]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302949.4]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302949.4]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302949.4]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302949.4]
  wire  AsyncResetRegVec_w1_i0_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302978.4]
  wire  AsyncResetRegVec_w1_i0_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302978.4]
  wire  AsyncResetRegVec_w1_i0_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302978.4]
  wire  AsyncResetRegVec_w1_i0_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302978.4]
  wire  AsyncResetRegVec_w1_i0_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302978.4]
  wire  _T_86; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302876.4]
  wire  source_ready; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302874.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302875.4 AsyncQueue.scala 164:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302964.4]
  wire  _T_87; // @[AsyncQueue.scala 130:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302877.4]
  wire [3:0] _GEN_24; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302885.4]
  wire [3:0] _T_91; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302886.4]
  wire [3:0] _T_92; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302887.4]
  wire [2:0] _T_93; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302889.4]
  wire [3:0] _GEN_25; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302890.4]
  wire [3:0] ridx; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302890.4]
  wire [3:0] widx; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302896.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302898.4]
  wire  _T_95; // @[AsyncQueue.scala 132:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302899.4]
  wire  valid; // @[AsyncQueue.scala 132:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302900.4]
  wire [2:0] _T_96; // @[AsyncQueue.scala 138:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302901.4]
  wire  _T_97; // @[AsyncQueue.scala 138:62:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302902.4]
  wire [2:0] _GEN_26; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302903.4]
  wire [2:0] _T_98; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302903.4]
  wire [2:0] index; // @[AsyncQueue.scala 138:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302904.4]
  wire [63:0] _GEN_3; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [7:0] _GEN_4; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire  _GEN_5; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [63:0] _GEN_6; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [7:0] _GEN_7; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire  _GEN_8; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [63:0] _GEN_9; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [7:0] _GEN_10; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire  _GEN_11; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [63:0] _GEN_12; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [7:0] _GEN_13; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire  _GEN_14; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [63:0] _GEN_15; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [7:0] _GEN_16; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire  _GEN_17; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [63:0] _GEN_18; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [7:0] _GEN_19; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire  _GEN_20; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [63:0] _GEN_21; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [7:0] _GEN_22; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire  _GEN_23; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [63:0] deq_bits_nxt_data; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [7:0] deq_bits_nxt_strb; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire  deq_bits_nxt_last; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  wire [71:0] _T_100; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302910.4]
  wire [72:0] _T_105; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302915.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302917.4]
  wire  valid_reg_1; // @[AsyncQueue.scala 147:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302933.4]
  wire  _T_111; // @[AsyncQueue.scala 157:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302953.4]
  AsyncResetRegVec_w4_i0 ridx_bin ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302879.4]
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_gray ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302891.4]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  SynchronizerShiftReg_w73_d1 deq_bits_reg ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302906.4]
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q)
  );
  AsyncResetRegVec_w1_i0 valid_reg ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302927.4]
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_w4_i0 ridx_gray ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302936.4]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302943.4]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302946.4]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302949.4]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302978.4]
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q),
    .io_en(AsyncResetRegVec_w1_i0_io_en)
  );
  assign _T_86 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302876.4]
  assign source_ready = AsyncValidSync_2_io_out; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302874.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302875.4 AsyncQueue.scala 164:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302964.4]
  assign _T_87 = source_ready == 1'h0; // @[AsyncQueue.scala 130:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302877.4]
  assign _GEN_24 = {{3'd0}, _T_86}; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302885.4]
  assign _T_91 = ridx_bin_io_q + _GEN_24; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302886.4]
  assign _T_92 = _T_87 ? 4'h0 : _T_91; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302887.4]
  assign _T_93 = _T_92[3:1]; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302889.4]
  assign _GEN_25 = {{1'd0}, _T_93}; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302890.4]
  assign ridx = _T_92 ^ _GEN_25; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302890.4]
  assign widx = widx_gray_io_q; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302896.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302898.4]
  assign _T_95 = ridx != widx; // @[AsyncQueue.scala 132:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302899.4]
  assign valid = source_ready & _T_95; // @[AsyncQueue.scala 132:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302900.4]
  assign _T_96 = ridx[2:0]; // @[AsyncQueue.scala 138:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302901.4]
  assign _T_97 = ridx[3]; // @[AsyncQueue.scala 138:62:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302902.4]
  assign _GEN_26 = {{2'd0}, _T_97}; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302903.4]
  assign _T_98 = _GEN_26 << 2; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302903.4]
  assign index = _T_96 ^ _T_98; // @[AsyncQueue.scala 138:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302904.4]
  assign _GEN_3 = 3'h1 == index ? io_async_mem_1_data : io_async_mem_0_data; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_4 = 3'h1 == index ? io_async_mem_1_strb : io_async_mem_0_strb; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_5 = 3'h1 == index ? io_async_mem_1_last : io_async_mem_0_last; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_6 = 3'h2 == index ? io_async_mem_2_data : _GEN_3; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_7 = 3'h2 == index ? io_async_mem_2_strb : _GEN_4; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_8 = 3'h2 == index ? io_async_mem_2_last : _GEN_5; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_9 = 3'h3 == index ? io_async_mem_3_data : _GEN_6; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_10 = 3'h3 == index ? io_async_mem_3_strb : _GEN_7; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_11 = 3'h3 == index ? io_async_mem_3_last : _GEN_8; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_12 = 3'h4 == index ? io_async_mem_4_data : _GEN_9; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_13 = 3'h4 == index ? io_async_mem_4_strb : _GEN_10; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_14 = 3'h4 == index ? io_async_mem_4_last : _GEN_11; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_15 = 3'h5 == index ? io_async_mem_5_data : _GEN_12; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_16 = 3'h5 == index ? io_async_mem_5_strb : _GEN_13; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_17 = 3'h5 == index ? io_async_mem_5_last : _GEN_14; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_18 = 3'h6 == index ? io_async_mem_6_data : _GEN_15; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_19 = 3'h6 == index ? io_async_mem_6_strb : _GEN_16; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_20 = 3'h6 == index ? io_async_mem_6_last : _GEN_17; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_21 = 3'h7 == index ? io_async_mem_7_data : _GEN_18; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_22 = 3'h7 == index ? io_async_mem_7_strb : _GEN_19; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _GEN_23 = 3'h7 == index ? io_async_mem_7_last : _GEN_20; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign deq_bits_nxt_data = valid ? _GEN_21 : io_deq_bits_data; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign deq_bits_nxt_strb = valid ? _GEN_22 : io_deq_bits_strb; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign deq_bits_nxt_last = valid ? _GEN_23 : io_deq_bits_last; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302905.4]
  assign _T_100 = {deq_bits_nxt_data,deq_bits_nxt_strb}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302910.4]
  assign _T_105 = deq_bits_reg_io_q; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302915.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302917.4]
  assign valid_reg_1 = valid_reg_io_q; // @[AsyncQueue.scala 147:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302933.4]
  assign _T_111 = io_async_safe_source_reset_n == 1'h0; // @[AsyncQueue.scala 157:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302953.4]
  assign io_deq_valid = valid_reg_1 & source_ready; // @[AsyncQueue.scala 148:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302935.4]
  assign io_deq_bits_data = _T_105[72:9]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302926.4]
  assign io_deq_bits_strb = _T_105[8:1]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302925.4]
  assign io_deq_bits_last = _T_105[0]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302924.4]
  assign io_async_ridx = ridx_gray_io_q; // @[AsyncQueue.scala 151:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302942.4]
  assign io_async_safe_ridx_valid = AsyncValidSync_io_out; // @[AsyncQueue.scala 161:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302961.4]
  assign io_async_safe_sink_reset_n = reset == 1'h0; // @[AsyncQueue.scala 165:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302967.4]
  assign ridx_bin_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302881.4]
  assign ridx_bin_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302882.4]
  assign ridx_bin_io_d = _T_87 ? 4'h0 : _T_91; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302883.4]
  assign ridx_bin_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302884.4]
  assign widx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302893.4]
  assign widx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302894.4]
  assign widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302895.4]
  assign deq_bits_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302908.4]
  assign deq_bits_reg_io_d = {_T_100,deq_bits_nxt_last}; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302912.4]
  assign valid_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302929.4]
  assign valid_reg_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302930.4]
  assign valid_reg_io_d = source_ready & _T_95; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302931.4]
  assign valid_reg_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302932.4]
  assign ridx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302938.4]
  assign ridx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302939.4]
  assign ridx_gray_io_d = _T_92 ^ _GEN_25; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302940.4]
  assign ridx_gray_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302941.4]
  assign AsyncValidSync_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302944.4]
  assign AsyncValidSync_reset = reset | _T_111; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302945.4 AsyncQueue.scala 157:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302955.4]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 160:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302960.4]
  assign AsyncValidSync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302947.4]
  assign AsyncValidSync_1_reset = reset | _T_111; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302948.4 AsyncQueue.scala 158:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302959.4]
  assign AsyncValidSync_1_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 162:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302962.4]
  assign AsyncValidSync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302950.4]
  assign AsyncValidSync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302951.4]
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 163:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302963.4]
  assign AsyncResetRegVec_w1_i0_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302980.4]
  assign AsyncResetRegVec_w1_i0_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302981.4]
  assign AsyncResetRegVec_w1_i0_io_d = io_async_widx == io_async_ridx; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302982.4]
  assign AsyncResetRegVec_w1_i0_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@302983.4]
endmodule
module AsyncQueueSource_3( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303900.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303901.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303902.4]
  output        io_enq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  input         io_enq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  input  [3:0]  io_enq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  input  [63:0] io_enq_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  input  [1:0]  io_enq_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  input         io_enq_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [63:0] io_async_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [1:0]  io_async_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [63:0] io_async_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [1:0]  io_async_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [63:0] io_async_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [1:0]  io_async_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [63:0] io_async_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [1:0]  io_async_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [63:0] io_async_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [1:0]  io_async_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [63:0] io_async_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [1:0]  io_async_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [63:0] io_async_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [1:0]  io_async_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [63:0] io_async_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [1:0]  io_async_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  input  [3:0]  io_async_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output [3:0]  io_async_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  input         io_async_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  output        io_async_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
  input         io_async_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303903.4]
);
  wire  widx_bin_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303911.4]
  wire  widx_bin_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303911.4]
  wire [3:0] widx_bin_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303911.4]
  wire [3:0] widx_bin_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303911.4]
  wire  widx_bin_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303911.4]
  wire  ridx_gray_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303923.4]
  wire  ridx_gray_reset; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303923.4]
  wire [3:0] ridx_gray_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303923.4]
  wire [3:0] ridx_gray_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303923.4]
  wire  ready_reg_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303945.4]
  wire  ready_reg_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303945.4]
  wire  ready_reg_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303945.4]
  wire  ready_reg_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303945.4]
  wire  ready_reg_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303945.4]
  wire  widx_gray_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303954.4]
  wire  widx_gray_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303954.4]
  wire [3:0] widx_gray_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303954.4]
  wire [3:0] widx_gray_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303954.4]
  wire  widx_gray_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303954.4]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303993.4]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303993.4]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303993.4]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303993.4]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303996.4]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303996.4]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303996.4]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303996.4]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303999.4]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303999.4]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303999.4]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303999.4]
  reg [3:0] mem_0_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_0;
  reg [63:0] mem_0_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [63:0] _RAND_1;
  reg [1:0] mem_0_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_2;
  reg  mem_0_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_3;
  reg [3:0] mem_1_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_4;
  reg [63:0] mem_1_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [63:0] _RAND_5;
  reg [1:0] mem_1_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_6;
  reg  mem_1_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_7;
  reg [3:0] mem_2_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_8;
  reg [63:0] mem_2_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [63:0] _RAND_9;
  reg [1:0] mem_2_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_10;
  reg  mem_2_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_11;
  reg [3:0] mem_3_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_12;
  reg [63:0] mem_3_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [63:0] _RAND_13;
  reg [1:0] mem_3_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_14;
  reg  mem_3_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_15;
  reg [3:0] mem_4_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_16;
  reg [63:0] mem_4_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [63:0] _RAND_17;
  reg [1:0] mem_4_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_18;
  reg  mem_4_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_19;
  reg [3:0] mem_5_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_20;
  reg [63:0] mem_5_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [63:0] _RAND_21;
  reg [1:0] mem_5_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_22;
  reg  mem_5_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_23;
  reg [3:0] mem_6_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_24;
  reg [63:0] mem_6_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [63:0] _RAND_25;
  reg [1:0] mem_6_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_26;
  reg  mem_6_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_27;
  reg [3:0] mem_7_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_28;
  reg [63:0] mem_7_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [63:0] _RAND_29;
  reg [1:0] mem_7_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_30;
  reg  mem_7_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303907.4]
  reg [31:0] _RAND_31;
  wire  _T_64; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303908.4]
  wire  sink_ready; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303905.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303906.4 AsyncQueue.scala 106:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304014.4]
  wire  _T_65; // @[AsyncQueue.scala 77:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303909.4]
  wire [3:0] _GEN_64; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303917.4]
  wire [3:0] _T_69; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303918.4]
  wire [3:0] _T_70; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303919.4]
  wire [2:0] _T_71; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303921.4]
  wire [3:0] _GEN_65; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303922.4]
  wire [3:0] widx; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303922.4]
  wire [3:0] ridx; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303928.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303930.4]
  wire [3:0] _T_73; // @[AsyncQueue.scala 79:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303931.4]
  wire  _T_74; // @[AsyncQueue.scala 79:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303932.4]
  wire [2:0] _T_75; // @[AsyncQueue.scala 81:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303934.4]
  wire  _T_76; // @[AsyncQueue.scala 81:80:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303935.4]
  wire [2:0] _GEN_66; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303936.4]
  wire [2:0] _T_77; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303936.4]
  wire [2:0] index; // @[AsyncQueue.scala 81:64:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303937.4]
  wire  ready_reg_1; // @[AsyncQueue.scala 84:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303951.4]
  wire  _T_82; // @[AsyncQueue.scala 99:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304003.4]
  AsyncResetRegVec_w4_i0 widx_bin ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303911.4]
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_gray ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303923.4]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  AsyncResetRegVec_w1_i0 ready_reg ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303945.4]
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_w4_i0 widx_gray ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303954.4]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303993.4]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303996.4]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303999.4]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign _T_64 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303908.4]
  assign sink_ready = AsyncValidSync_2_io_out; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303905.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303906.4 AsyncQueue.scala 106:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304014.4]
  assign _T_65 = sink_ready == 1'h0; // @[AsyncQueue.scala 77:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303909.4]
  assign _GEN_64 = {{3'd0}, _T_64}; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303917.4]
  assign _T_69 = widx_bin_io_q + _GEN_64; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303918.4]
  assign _T_70 = _T_65 ? 4'h0 : _T_69; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303919.4]
  assign _T_71 = _T_70[3:1]; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303921.4]
  assign _GEN_65 = {{1'd0}, _T_71}; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303922.4]
  assign widx = _T_70 ^ _GEN_65; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303922.4]
  assign ridx = ridx_gray_io_q; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303928.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303930.4]
  assign _T_73 = ridx ^ 4'hc; // @[AsyncQueue.scala 79:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303931.4]
  assign _T_74 = widx != _T_73; // @[AsyncQueue.scala 79:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303932.4]
  assign _T_75 = io_async_widx[2:0]; // @[AsyncQueue.scala 81:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303934.4]
  assign _T_76 = io_async_widx[3]; // @[AsyncQueue.scala 81:80:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303935.4]
  assign _GEN_66 = {{2'd0}, _T_76}; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303936.4]
  assign _T_77 = _GEN_66 << 2; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303936.4]
  assign index = _T_75 ^ _T_77; // @[AsyncQueue.scala 81:64:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303937.4]
  assign ready_reg_1 = ready_reg_io_q; // @[AsyncQueue.scala 84:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303951.4]
  assign _T_82 = io_async_safe_sink_reset_n == 1'h0; // @[AsyncQueue.scala 99:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304003.4]
  assign io_enq_ready = ready_reg_1 & sink_ready; // @[AsyncQueue.scala 85:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303953.4]
  assign io_async_mem_0_id = mem_0_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303964.4]
  assign io_async_mem_0_data = mem_0_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303963.4]
  assign io_async_mem_0_resp = mem_0_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303962.4]
  assign io_async_mem_0_last = mem_0_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303961.4]
  assign io_async_mem_1_id = mem_1_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303968.4]
  assign io_async_mem_1_data = mem_1_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303967.4]
  assign io_async_mem_1_resp = mem_1_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303966.4]
  assign io_async_mem_1_last = mem_1_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303965.4]
  assign io_async_mem_2_id = mem_2_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303972.4]
  assign io_async_mem_2_data = mem_2_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303971.4]
  assign io_async_mem_2_resp = mem_2_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303970.4]
  assign io_async_mem_2_last = mem_2_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303969.4]
  assign io_async_mem_3_id = mem_3_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303976.4]
  assign io_async_mem_3_data = mem_3_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303975.4]
  assign io_async_mem_3_resp = mem_3_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303974.4]
  assign io_async_mem_3_last = mem_3_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303973.4]
  assign io_async_mem_4_id = mem_4_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303980.4]
  assign io_async_mem_4_data = mem_4_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303979.4]
  assign io_async_mem_4_resp = mem_4_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303978.4]
  assign io_async_mem_4_last = mem_4_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303977.4]
  assign io_async_mem_5_id = mem_5_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303984.4]
  assign io_async_mem_5_data = mem_5_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303983.4]
  assign io_async_mem_5_resp = mem_5_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303982.4]
  assign io_async_mem_5_last = mem_5_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303981.4]
  assign io_async_mem_6_id = mem_6_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303988.4]
  assign io_async_mem_6_data = mem_6_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303987.4]
  assign io_async_mem_6_resp = mem_6_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303986.4]
  assign io_async_mem_6_last = mem_6_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303985.4]
  assign io_async_mem_7_id = mem_7_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303992.4]
  assign io_async_mem_7_data = mem_7_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303991.4]
  assign io_async_mem_7_resp = mem_7_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303990.4]
  assign io_async_mem_7_last = mem_7_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303989.4]
  assign io_async_widx = widx_gray_io_q; // @[AsyncQueue.scala 88:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303960.4]
  assign io_async_safe_widx_valid = AsyncValidSync_io_out; // @[AsyncQueue.scala 103:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304011.4]
  assign io_async_safe_source_reset_n = reset == 1'h0; // @[AsyncQueue.scala 107:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304017.4]
  assign widx_bin_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303913.4]
  assign widx_bin_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303914.4]
  assign widx_bin_io_d = _T_65 ? 4'h0 : _T_69; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303915.4]
  assign widx_bin_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303916.4]
  assign ridx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303925.4]
  assign ridx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303926.4]
  assign ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303927.4]
  assign ready_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303947.4]
  assign ready_reg_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303948.4]
  assign ready_reg_io_d = sink_ready & _T_74; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303949.4]
  assign ready_reg_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303950.4]
  assign widx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303956.4]
  assign widx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303957.4]
  assign widx_gray_io_d = _T_70 ^ _GEN_65; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303958.4]
  assign widx_gray_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303959.4]
  assign AsyncValidSync_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303994.4]
  assign AsyncValidSync_reset = reset | _T_82; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303995.4 AsyncQueue.scala 99:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304005.4]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 102:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304010.4]
  assign AsyncValidSync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303997.4]
  assign AsyncValidSync_1_reset = reset | _T_82; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@303998.4 AsyncQueue.scala 100:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304009.4]
  assign AsyncValidSync_1_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 104:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304012.4]
  assign AsyncValidSync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304000.4]
  assign AsyncValidSync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304001.4]
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 105:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304013.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_id = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  mem_0_data = _RAND_1[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_0_resp = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_0_last = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_1_id = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  mem_1_data = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_1_resp = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_1_last = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_2_id = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  mem_2_data = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_2_resp = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_2_last = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mem_3_id = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  mem_3_data = _RAND_13[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mem_3_resp = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mem_3_last = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  mem_4_id = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  mem_4_data = _RAND_17[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  mem_4_resp = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  mem_4_last = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  mem_5_id = _RAND_20[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  mem_5_data = _RAND_21[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_5_resp = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_5_last = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mem_6_id = _RAND_24[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  mem_6_data = _RAND_25[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_6_resp = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_6_last = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_7_id = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  mem_7_data = _RAND_29[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_7_resp = _RAND_30[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_7_last = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_last <= io_enq_bits_last;
      end
    end
  end
endmodule
module AsyncQueueSource_4( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304934.2]
  input        clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304935.4]
  input        reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304936.4]
  output       io_enq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  input        io_enq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  input  [3:0] io_enq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  input  [1:0] io_enq_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [1:0] io_async_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [1:0] io_async_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [1:0] io_async_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [1:0] io_async_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [1:0] io_async_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [1:0] io_async_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [1:0] io_async_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [1:0] io_async_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  input  [3:0] io_async_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output [3:0] io_async_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  input        io_async_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output       io_async_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  output       io_async_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
  input        io_async_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304937.4]
);
  wire  widx_bin_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304945.4]
  wire  widx_bin_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304945.4]
  wire [3:0] widx_bin_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304945.4]
  wire [3:0] widx_bin_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304945.4]
  wire  widx_bin_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304945.4]
  wire  ridx_gray_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304957.4]
  wire  ridx_gray_reset; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304957.4]
  wire [3:0] ridx_gray_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304957.4]
  wire [3:0] ridx_gray_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304957.4]
  wire  ready_reg_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304977.4]
  wire  ready_reg_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304977.4]
  wire  ready_reg_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304977.4]
  wire  ready_reg_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304977.4]
  wire  ready_reg_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304977.4]
  wire  widx_gray_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304986.4]
  wire  widx_gray_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304986.4]
  wire [3:0] widx_gray_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304986.4]
  wire [3:0] widx_gray_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304986.4]
  wire  widx_gray_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304986.4]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305009.4]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305009.4]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305009.4]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305009.4]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305012.4]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305012.4]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305012.4]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305012.4]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305015.4]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305015.4]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305015.4]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305015.4]
  reg [3:0] mem_0_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_0;
  reg [1:0] mem_0_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_1;
  reg [3:0] mem_1_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_2;
  reg [1:0] mem_1_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_3;
  reg [3:0] mem_2_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_4;
  reg [1:0] mem_2_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_5;
  reg [3:0] mem_3_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_6;
  reg [1:0] mem_3_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_7;
  reg [3:0] mem_4_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_8;
  reg [1:0] mem_4_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_9;
  reg [3:0] mem_5_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_10;
  reg [1:0] mem_5_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_11;
  reg [3:0] mem_6_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_12;
  reg [1:0] mem_6_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_13;
  reg [3:0] mem_7_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_14;
  reg [1:0] mem_7_resp; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304941.4]
  reg [31:0] _RAND_15;
  wire  _T_64; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304942.4]
  wire  sink_ready; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304939.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304940.4 AsyncQueue.scala 106:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305030.4]
  wire  _T_65; // @[AsyncQueue.scala 77:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304943.4]
  wire [3:0] _GEN_32; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304951.4]
  wire [3:0] _T_69; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304952.4]
  wire [3:0] _T_70; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304953.4]
  wire [2:0] _T_71; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304955.4]
  wire [3:0] _GEN_33; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304956.4]
  wire [3:0] widx; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304956.4]
  wire [3:0] ridx; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304962.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304964.4]
  wire [3:0] _T_73; // @[AsyncQueue.scala 79:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304965.4]
  wire  _T_74; // @[AsyncQueue.scala 79:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304966.4]
  wire [2:0] _T_75; // @[AsyncQueue.scala 81:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304968.4]
  wire  _T_76; // @[AsyncQueue.scala 81:80:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304969.4]
  wire [2:0] _GEN_34; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304970.4]
  wire [2:0] _T_77; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304970.4]
  wire [2:0] index; // @[AsyncQueue.scala 81:64:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304971.4]
  wire  ready_reg_1; // @[AsyncQueue.scala 84:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304983.4]
  wire  _T_82; // @[AsyncQueue.scala 99:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305019.4]
  AsyncResetRegVec_w4_i0 widx_bin ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304945.4]
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_gray ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304957.4]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  AsyncResetRegVec_w1_i0 ready_reg ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304977.4]
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_w4_i0 widx_gray ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304986.4]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305009.4]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305012.4]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305015.4]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign _T_64 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304942.4]
  assign sink_ready = AsyncValidSync_2_io_out; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304939.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304940.4 AsyncQueue.scala 106:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305030.4]
  assign _T_65 = sink_ready == 1'h0; // @[AsyncQueue.scala 77:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304943.4]
  assign _GEN_32 = {{3'd0}, _T_64}; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304951.4]
  assign _T_69 = widx_bin_io_q + _GEN_32; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304952.4]
  assign _T_70 = _T_65 ? 4'h0 : _T_69; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304953.4]
  assign _T_71 = _T_70[3:1]; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304955.4]
  assign _GEN_33 = {{1'd0}, _T_71}; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304956.4]
  assign widx = _T_70 ^ _GEN_33; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304956.4]
  assign ridx = ridx_gray_io_q; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304962.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304964.4]
  assign _T_73 = ridx ^ 4'hc; // @[AsyncQueue.scala 79:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304965.4]
  assign _T_74 = widx != _T_73; // @[AsyncQueue.scala 79:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304966.4]
  assign _T_75 = io_async_widx[2:0]; // @[AsyncQueue.scala 81:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304968.4]
  assign _T_76 = io_async_widx[3]; // @[AsyncQueue.scala 81:80:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304969.4]
  assign _GEN_34 = {{2'd0}, _T_76}; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304970.4]
  assign _T_77 = _GEN_34 << 2; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304970.4]
  assign index = _T_75 ^ _T_77; // @[AsyncQueue.scala 81:64:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304971.4]
  assign ready_reg_1 = ready_reg_io_q; // @[AsyncQueue.scala 84:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304983.4]
  assign _T_82 = io_async_safe_sink_reset_n == 1'h0; // @[AsyncQueue.scala 99:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305019.4]
  assign io_enq_ready = ready_reg_1 & sink_ready; // @[AsyncQueue.scala 85:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304985.4]
  assign io_async_mem_0_id = mem_0_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304994.4]
  assign io_async_mem_0_resp = mem_0_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304993.4]
  assign io_async_mem_1_id = mem_1_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304996.4]
  assign io_async_mem_1_resp = mem_1_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304995.4]
  assign io_async_mem_2_id = mem_2_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304998.4]
  assign io_async_mem_2_resp = mem_2_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304997.4]
  assign io_async_mem_3_id = mem_3_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305000.4]
  assign io_async_mem_3_resp = mem_3_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304999.4]
  assign io_async_mem_4_id = mem_4_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305002.4]
  assign io_async_mem_4_resp = mem_4_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305001.4]
  assign io_async_mem_5_id = mem_5_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305004.4]
  assign io_async_mem_5_resp = mem_5_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305003.4]
  assign io_async_mem_6_id = mem_6_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305006.4]
  assign io_async_mem_6_resp = mem_6_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305005.4]
  assign io_async_mem_7_id = mem_7_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305008.4]
  assign io_async_mem_7_resp = mem_7_resp; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305007.4]
  assign io_async_widx = widx_gray_io_q; // @[AsyncQueue.scala 88:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304992.4]
  assign io_async_safe_widx_valid = AsyncValidSync_io_out; // @[AsyncQueue.scala 103:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305027.4]
  assign io_async_safe_source_reset_n = reset == 1'h0; // @[AsyncQueue.scala 107:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305033.4]
  assign widx_bin_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304947.4]
  assign widx_bin_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304948.4]
  assign widx_bin_io_d = _T_65 ? 4'h0 : _T_69; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304949.4]
  assign widx_bin_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304950.4]
  assign ridx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304959.4]
  assign ridx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304960.4]
  assign ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304961.4]
  assign ready_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304979.4]
  assign ready_reg_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304980.4]
  assign ready_reg_io_d = sink_ready & _T_74; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304981.4]
  assign ready_reg_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304982.4]
  assign widx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304988.4]
  assign widx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304989.4]
  assign widx_gray_io_d = _T_70 ^ _GEN_33; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304990.4]
  assign widx_gray_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@304991.4]
  assign AsyncValidSync_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305010.4]
  assign AsyncValidSync_reset = reset | _T_82; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305011.4 AsyncQueue.scala 99:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305021.4]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 102:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305026.4]
  assign AsyncValidSync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305013.4]
  assign AsyncValidSync_1_reset = reset | _T_82; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305014.4 AsyncQueue.scala 100:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305025.4]
  assign AsyncValidSync_1_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 104:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305028.4]
  assign AsyncValidSync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305016.4]
  assign AsyncValidSync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305017.4]
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 105:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305029.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_id = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_0_resp = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_1_id = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_1_resp = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_2_id = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_2_resp = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_3_id = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_3_resp = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_4_id = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mem_4_resp = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_5_id = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_5_resp = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mem_6_id = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mem_6_resp = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mem_7_id = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mem_7_resp = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_resp <= io_enq_bits_resp;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_resp <= io_enq_bits_resp;
      end
    end
  end
endmodule
module AXI4AsyncCrossingSink( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305035.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305036.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305037.4]
  input  [3:0]  auto_in_aw_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_aw_mem_0_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_aw_mem_0_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_0_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_aw_mem_0_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_mem_0_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_0_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_0_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_0_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_aw_mem_1_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_aw_mem_1_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_1_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_aw_mem_1_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_mem_1_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_1_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_1_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_1_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_aw_mem_2_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_aw_mem_2_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_2_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_aw_mem_2_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_mem_2_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_2_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_2_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_2_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_aw_mem_3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_aw_mem_3_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_3_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_aw_mem_3_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_mem_3_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_3_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_3_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_3_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_aw_mem_4_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_aw_mem_4_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_4_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_aw_mem_4_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_mem_4_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_4_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_4_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_4_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_aw_mem_5_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_aw_mem_5_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_5_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_aw_mem_5_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_mem_5_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_5_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_5_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_5_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_aw_mem_6_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_aw_mem_6_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_6_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_aw_mem_6_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_mem_6_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_6_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_6_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_6_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_aw_mem_7_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_aw_mem_7_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_7_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_aw_mem_7_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_mem_7_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_7_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_aw_mem_7_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_mem_7_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_aw_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_aw_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_aw_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_aw_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_aw_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_in_w_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_w_mem_0_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_in_w_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_w_mem_1_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_in_w_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_w_mem_2_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_in_w_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_w_mem_3_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_in_w_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_w_mem_4_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_in_w_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_w_mem_5_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_in_w_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_w_mem_6_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_in_w_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_w_mem_7_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_w_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_w_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_w_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_w_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_w_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_b_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_b_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_b_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_b_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_b_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_b_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_b_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_b_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_b_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_b_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_b_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_b_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_b_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_b_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_ar_mem_0_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_ar_mem_0_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_0_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_ar_mem_0_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_mem_0_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_0_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_0_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_0_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_ar_mem_1_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_ar_mem_1_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_1_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_ar_mem_1_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_mem_1_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_1_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_1_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_1_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_ar_mem_2_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_ar_mem_2_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_2_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_ar_mem_2_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_mem_2_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_2_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_2_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_2_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_ar_mem_3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_ar_mem_3_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_3_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_ar_mem_3_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_mem_3_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_3_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_3_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_3_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_ar_mem_4_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_ar_mem_4_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_4_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_ar_mem_4_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_mem_4_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_4_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_4_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_4_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_ar_mem_5_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_ar_mem_5_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_5_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_ar_mem_5_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_mem_5_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_5_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_5_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_5_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_ar_mem_6_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_ar_mem_6_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_6_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_ar_mem_6_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_mem_6_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_6_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_6_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_6_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [31:0] auto_in_ar_mem_7_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [7:0]  auto_in_ar_mem_7_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_7_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_in_ar_mem_7_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_mem_7_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_7_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [2:0]  auto_in_ar_mem_7_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_mem_7_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_ar_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_ar_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_ar_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_ar_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_ar_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_in_r_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_r_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_in_r_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_r_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_in_r_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_r_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_in_r_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_r_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_in_r_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_r_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_in_r_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_r_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_in_r_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_r_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_in_r_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_in_r_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_in_r_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_in_r_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_r_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_in_r_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_in_r_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_out_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_out_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_out_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [31:0] auto_out_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [7:0]  auto_out_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [2:0]  auto_out_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_out_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_out_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_out_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [63:0] auto_out_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [7:0]  auto_out_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_out_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_out_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_out_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_out_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_out_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_out_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_out_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [31:0] auto_out_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [7:0]  auto_out_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [2:0]  auto_out_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_out_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  output        auto_out_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_out_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [3:0]  auto_out_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [63:0] auto_out_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
  input         auto_out_r_bits_last // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305038.4]
);
  wire  AsyncQueueSink_clock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_reset; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_deq_ready; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_deq_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_deq_bits_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_deq_bits_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_deq_bits_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_deq_bits_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_deq_bits_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_deq_bits_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_deq_bits_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_deq_bits_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_deq_bits_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_0_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_async_mem_0_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_async_mem_0_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_0_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_async_mem_0_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_mem_0_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_0_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_0_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_0_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_1_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_async_mem_1_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_async_mem_1_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_1_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_async_mem_1_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_mem_1_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_1_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_1_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_1_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_2_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_async_mem_2_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_async_mem_2_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_2_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_async_mem_2_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_mem_2_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_2_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_2_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_2_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_3_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_async_mem_3_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_async_mem_3_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_3_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_async_mem_3_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_mem_3_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_3_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_3_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_3_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_4_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_async_mem_4_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_async_mem_4_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_4_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_async_mem_4_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_mem_4_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_4_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_4_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_4_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_5_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_async_mem_5_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_async_mem_5_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_5_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_async_mem_5_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_mem_5_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_5_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_5_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_5_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_6_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_async_mem_6_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_async_mem_6_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_6_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_async_mem_6_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_mem_6_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_6_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_6_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_6_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_7_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [31:0] AsyncQueueSink_io_async_mem_7_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [7:0] AsyncQueueSink_io_async_mem_7_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_7_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [1:0] AsyncQueueSink_io_async_mem_7_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_mem_7_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_7_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [2:0] AsyncQueueSink_io_async_mem_7_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_mem_7_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_ridx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire [3:0] AsyncQueueSink_io_async_widx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_safe_widx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
  wire  AsyncQueueSink_1_clock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_reset; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_deq_ready; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_deq_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_deq_bits_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_deq_bits_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_deq_bits_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_deq_bits_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_deq_bits_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_deq_bits_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_deq_bits_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_deq_bits_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_deq_bits_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_0_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_async_mem_0_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_async_mem_0_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_0_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_0_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_mem_0_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_0_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_0_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_0_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_1_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_async_mem_1_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_async_mem_1_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_1_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_1_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_mem_1_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_1_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_1_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_1_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_2_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_async_mem_2_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_async_mem_2_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_2_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_2_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_mem_2_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_2_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_2_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_2_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_3_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_async_mem_3_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_async_mem_3_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_3_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_3_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_mem_3_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_3_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_3_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_3_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_4_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_async_mem_4_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_async_mem_4_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_4_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_4_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_mem_4_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_4_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_4_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_4_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_5_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_async_mem_5_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_async_mem_5_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_5_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_5_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_mem_5_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_5_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_5_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_5_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_6_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_async_mem_6_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_async_mem_6_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_6_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_6_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_mem_6_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_6_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_6_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_6_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_7_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [31:0] AsyncQueueSink_1_io_async_mem_7_addr; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [7:0] AsyncQueueSink_1_io_async_mem_7_len; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_7_size; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_7_burst; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_mem_7_lock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_7_cache; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [2:0] AsyncQueueSink_1_io_async_mem_7_prot; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_7_qos; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_ridx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire [3:0] AsyncQueueSink_1_io_async_widx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_safe_ridx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_safe_widx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_safe_source_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_1_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
  wire  AsyncQueueSink_2_clock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_reset; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_deq_ready; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_deq_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_deq_bits_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_deq_bits_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_deq_bits_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_async_mem_0_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_async_mem_0_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_mem_0_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_async_mem_1_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_async_mem_1_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_mem_1_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_async_mem_2_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_async_mem_2_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_mem_2_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_async_mem_3_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_async_mem_3_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_mem_3_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_async_mem_4_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_async_mem_4_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_mem_4_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_async_mem_5_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_async_mem_5_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_mem_5_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_async_mem_6_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_async_mem_6_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_mem_6_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [63:0] AsyncQueueSink_2_io_async_mem_7_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [7:0] AsyncQueueSink_2_io_async_mem_7_strb; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_mem_7_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [3:0] AsyncQueueSink_2_io_async_ridx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire [3:0] AsyncQueueSink_2_io_async_widx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_safe_ridx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_safe_widx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_safe_source_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSink_2_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
  wire  AsyncQueueSource_clock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_reset; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_enq_ready; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_enq_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_enq_bits_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_enq_bits_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_enq_bits_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_enq_bits_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_mem_0_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_async_mem_0_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_async_mem_0_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_mem_0_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_mem_1_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_async_mem_1_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_async_mem_1_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_mem_1_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_mem_2_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_async_mem_2_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_async_mem_2_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_mem_2_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_mem_3_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_async_mem_3_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_async_mem_3_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_mem_3_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_mem_4_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_async_mem_4_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_async_mem_4_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_mem_4_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_mem_5_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_async_mem_5_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_async_mem_5_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_mem_5_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_mem_6_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_async_mem_6_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_async_mem_6_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_mem_6_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_mem_7_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [63:0] AsyncQueueSource_io_async_mem_7_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [1:0] AsyncQueueSource_io_async_mem_7_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_mem_7_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_ridx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire [3:0] AsyncQueueSource_io_async_widx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_safe_ridx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_safe_widx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_safe_source_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
  wire  AsyncQueueSource_1_clock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire  AsyncQueueSource_1_reset; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire  AsyncQueueSource_1_io_enq_ready; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire  AsyncQueueSource_1_io_enq_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_enq_bits_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_enq_bits_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_0_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_0_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_1_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_1_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_2_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_2_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_3_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_3_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_4_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_4_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_5_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_5_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_6_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_6_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_7_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_7_resp; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_ridx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire [3:0] AsyncQueueSource_1_io_async_widx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire  AsyncQueueSource_1_io_async_safe_ridx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire  AsyncQueueSource_1_io_async_safe_widx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire  AsyncQueueSource_1_io_async_safe_source_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  wire  AsyncQueueSource_1_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
  AsyncQueueSink_3 AsyncQueueSink ( // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305049.4]
    .clock(AsyncQueueSink_clock),
    .reset(AsyncQueueSink_reset),
    .io_deq_ready(AsyncQueueSink_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_io_deq_valid),
    .io_deq_bits_id(AsyncQueueSink_io_deq_bits_id),
    .io_deq_bits_addr(AsyncQueueSink_io_deq_bits_addr),
    .io_deq_bits_len(AsyncQueueSink_io_deq_bits_len),
    .io_deq_bits_size(AsyncQueueSink_io_deq_bits_size),
    .io_deq_bits_burst(AsyncQueueSink_io_deq_bits_burst),
    .io_deq_bits_lock(AsyncQueueSink_io_deq_bits_lock),
    .io_deq_bits_cache(AsyncQueueSink_io_deq_bits_cache),
    .io_deq_bits_prot(AsyncQueueSink_io_deq_bits_prot),
    .io_deq_bits_qos(AsyncQueueSink_io_deq_bits_qos),
    .io_async_mem_0_id(AsyncQueueSink_io_async_mem_0_id),
    .io_async_mem_0_addr(AsyncQueueSink_io_async_mem_0_addr),
    .io_async_mem_0_len(AsyncQueueSink_io_async_mem_0_len),
    .io_async_mem_0_size(AsyncQueueSink_io_async_mem_0_size),
    .io_async_mem_0_burst(AsyncQueueSink_io_async_mem_0_burst),
    .io_async_mem_0_lock(AsyncQueueSink_io_async_mem_0_lock),
    .io_async_mem_0_cache(AsyncQueueSink_io_async_mem_0_cache),
    .io_async_mem_0_prot(AsyncQueueSink_io_async_mem_0_prot),
    .io_async_mem_0_qos(AsyncQueueSink_io_async_mem_0_qos),
    .io_async_mem_1_id(AsyncQueueSink_io_async_mem_1_id),
    .io_async_mem_1_addr(AsyncQueueSink_io_async_mem_1_addr),
    .io_async_mem_1_len(AsyncQueueSink_io_async_mem_1_len),
    .io_async_mem_1_size(AsyncQueueSink_io_async_mem_1_size),
    .io_async_mem_1_burst(AsyncQueueSink_io_async_mem_1_burst),
    .io_async_mem_1_lock(AsyncQueueSink_io_async_mem_1_lock),
    .io_async_mem_1_cache(AsyncQueueSink_io_async_mem_1_cache),
    .io_async_mem_1_prot(AsyncQueueSink_io_async_mem_1_prot),
    .io_async_mem_1_qos(AsyncQueueSink_io_async_mem_1_qos),
    .io_async_mem_2_id(AsyncQueueSink_io_async_mem_2_id),
    .io_async_mem_2_addr(AsyncQueueSink_io_async_mem_2_addr),
    .io_async_mem_2_len(AsyncQueueSink_io_async_mem_2_len),
    .io_async_mem_2_size(AsyncQueueSink_io_async_mem_2_size),
    .io_async_mem_2_burst(AsyncQueueSink_io_async_mem_2_burst),
    .io_async_mem_2_lock(AsyncQueueSink_io_async_mem_2_lock),
    .io_async_mem_2_cache(AsyncQueueSink_io_async_mem_2_cache),
    .io_async_mem_2_prot(AsyncQueueSink_io_async_mem_2_prot),
    .io_async_mem_2_qos(AsyncQueueSink_io_async_mem_2_qos),
    .io_async_mem_3_id(AsyncQueueSink_io_async_mem_3_id),
    .io_async_mem_3_addr(AsyncQueueSink_io_async_mem_3_addr),
    .io_async_mem_3_len(AsyncQueueSink_io_async_mem_3_len),
    .io_async_mem_3_size(AsyncQueueSink_io_async_mem_3_size),
    .io_async_mem_3_burst(AsyncQueueSink_io_async_mem_3_burst),
    .io_async_mem_3_lock(AsyncQueueSink_io_async_mem_3_lock),
    .io_async_mem_3_cache(AsyncQueueSink_io_async_mem_3_cache),
    .io_async_mem_3_prot(AsyncQueueSink_io_async_mem_3_prot),
    .io_async_mem_3_qos(AsyncQueueSink_io_async_mem_3_qos),
    .io_async_mem_4_id(AsyncQueueSink_io_async_mem_4_id),
    .io_async_mem_4_addr(AsyncQueueSink_io_async_mem_4_addr),
    .io_async_mem_4_len(AsyncQueueSink_io_async_mem_4_len),
    .io_async_mem_4_size(AsyncQueueSink_io_async_mem_4_size),
    .io_async_mem_4_burst(AsyncQueueSink_io_async_mem_4_burst),
    .io_async_mem_4_lock(AsyncQueueSink_io_async_mem_4_lock),
    .io_async_mem_4_cache(AsyncQueueSink_io_async_mem_4_cache),
    .io_async_mem_4_prot(AsyncQueueSink_io_async_mem_4_prot),
    .io_async_mem_4_qos(AsyncQueueSink_io_async_mem_4_qos),
    .io_async_mem_5_id(AsyncQueueSink_io_async_mem_5_id),
    .io_async_mem_5_addr(AsyncQueueSink_io_async_mem_5_addr),
    .io_async_mem_5_len(AsyncQueueSink_io_async_mem_5_len),
    .io_async_mem_5_size(AsyncQueueSink_io_async_mem_5_size),
    .io_async_mem_5_burst(AsyncQueueSink_io_async_mem_5_burst),
    .io_async_mem_5_lock(AsyncQueueSink_io_async_mem_5_lock),
    .io_async_mem_5_cache(AsyncQueueSink_io_async_mem_5_cache),
    .io_async_mem_5_prot(AsyncQueueSink_io_async_mem_5_prot),
    .io_async_mem_5_qos(AsyncQueueSink_io_async_mem_5_qos),
    .io_async_mem_6_id(AsyncQueueSink_io_async_mem_6_id),
    .io_async_mem_6_addr(AsyncQueueSink_io_async_mem_6_addr),
    .io_async_mem_6_len(AsyncQueueSink_io_async_mem_6_len),
    .io_async_mem_6_size(AsyncQueueSink_io_async_mem_6_size),
    .io_async_mem_6_burst(AsyncQueueSink_io_async_mem_6_burst),
    .io_async_mem_6_lock(AsyncQueueSink_io_async_mem_6_lock),
    .io_async_mem_6_cache(AsyncQueueSink_io_async_mem_6_cache),
    .io_async_mem_6_prot(AsyncQueueSink_io_async_mem_6_prot),
    .io_async_mem_6_qos(AsyncQueueSink_io_async_mem_6_qos),
    .io_async_mem_7_id(AsyncQueueSink_io_async_mem_7_id),
    .io_async_mem_7_addr(AsyncQueueSink_io_async_mem_7_addr),
    .io_async_mem_7_len(AsyncQueueSink_io_async_mem_7_len),
    .io_async_mem_7_size(AsyncQueueSink_io_async_mem_7_size),
    .io_async_mem_7_burst(AsyncQueueSink_io_async_mem_7_burst),
    .io_async_mem_7_lock(AsyncQueueSink_io_async_mem_7_lock),
    .io_async_mem_7_cache(AsyncQueueSink_io_async_mem_7_cache),
    .io_async_mem_7_prot(AsyncQueueSink_io_async_mem_7_prot),
    .io_async_mem_7_qos(AsyncQueueSink_io_async_mem_7_qos),
    .io_async_ridx(AsyncQueueSink_io_async_ridx),
    .io_async_widx(AsyncQueueSink_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink_3 AsyncQueueSink_1 ( // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305067.4]
    .clock(AsyncQueueSink_1_clock),
    .reset(AsyncQueueSink_1_reset),
    .io_deq_ready(AsyncQueueSink_1_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_1_io_deq_valid),
    .io_deq_bits_id(AsyncQueueSink_1_io_deq_bits_id),
    .io_deq_bits_addr(AsyncQueueSink_1_io_deq_bits_addr),
    .io_deq_bits_len(AsyncQueueSink_1_io_deq_bits_len),
    .io_deq_bits_size(AsyncQueueSink_1_io_deq_bits_size),
    .io_deq_bits_burst(AsyncQueueSink_1_io_deq_bits_burst),
    .io_deq_bits_lock(AsyncQueueSink_1_io_deq_bits_lock),
    .io_deq_bits_cache(AsyncQueueSink_1_io_deq_bits_cache),
    .io_deq_bits_prot(AsyncQueueSink_1_io_deq_bits_prot),
    .io_deq_bits_qos(AsyncQueueSink_1_io_deq_bits_qos),
    .io_async_mem_0_id(AsyncQueueSink_1_io_async_mem_0_id),
    .io_async_mem_0_addr(AsyncQueueSink_1_io_async_mem_0_addr),
    .io_async_mem_0_len(AsyncQueueSink_1_io_async_mem_0_len),
    .io_async_mem_0_size(AsyncQueueSink_1_io_async_mem_0_size),
    .io_async_mem_0_burst(AsyncQueueSink_1_io_async_mem_0_burst),
    .io_async_mem_0_lock(AsyncQueueSink_1_io_async_mem_0_lock),
    .io_async_mem_0_cache(AsyncQueueSink_1_io_async_mem_0_cache),
    .io_async_mem_0_prot(AsyncQueueSink_1_io_async_mem_0_prot),
    .io_async_mem_0_qos(AsyncQueueSink_1_io_async_mem_0_qos),
    .io_async_mem_1_id(AsyncQueueSink_1_io_async_mem_1_id),
    .io_async_mem_1_addr(AsyncQueueSink_1_io_async_mem_1_addr),
    .io_async_mem_1_len(AsyncQueueSink_1_io_async_mem_1_len),
    .io_async_mem_1_size(AsyncQueueSink_1_io_async_mem_1_size),
    .io_async_mem_1_burst(AsyncQueueSink_1_io_async_mem_1_burst),
    .io_async_mem_1_lock(AsyncQueueSink_1_io_async_mem_1_lock),
    .io_async_mem_1_cache(AsyncQueueSink_1_io_async_mem_1_cache),
    .io_async_mem_1_prot(AsyncQueueSink_1_io_async_mem_1_prot),
    .io_async_mem_1_qos(AsyncQueueSink_1_io_async_mem_1_qos),
    .io_async_mem_2_id(AsyncQueueSink_1_io_async_mem_2_id),
    .io_async_mem_2_addr(AsyncQueueSink_1_io_async_mem_2_addr),
    .io_async_mem_2_len(AsyncQueueSink_1_io_async_mem_2_len),
    .io_async_mem_2_size(AsyncQueueSink_1_io_async_mem_2_size),
    .io_async_mem_2_burst(AsyncQueueSink_1_io_async_mem_2_burst),
    .io_async_mem_2_lock(AsyncQueueSink_1_io_async_mem_2_lock),
    .io_async_mem_2_cache(AsyncQueueSink_1_io_async_mem_2_cache),
    .io_async_mem_2_prot(AsyncQueueSink_1_io_async_mem_2_prot),
    .io_async_mem_2_qos(AsyncQueueSink_1_io_async_mem_2_qos),
    .io_async_mem_3_id(AsyncQueueSink_1_io_async_mem_3_id),
    .io_async_mem_3_addr(AsyncQueueSink_1_io_async_mem_3_addr),
    .io_async_mem_3_len(AsyncQueueSink_1_io_async_mem_3_len),
    .io_async_mem_3_size(AsyncQueueSink_1_io_async_mem_3_size),
    .io_async_mem_3_burst(AsyncQueueSink_1_io_async_mem_3_burst),
    .io_async_mem_3_lock(AsyncQueueSink_1_io_async_mem_3_lock),
    .io_async_mem_3_cache(AsyncQueueSink_1_io_async_mem_3_cache),
    .io_async_mem_3_prot(AsyncQueueSink_1_io_async_mem_3_prot),
    .io_async_mem_3_qos(AsyncQueueSink_1_io_async_mem_3_qos),
    .io_async_mem_4_id(AsyncQueueSink_1_io_async_mem_4_id),
    .io_async_mem_4_addr(AsyncQueueSink_1_io_async_mem_4_addr),
    .io_async_mem_4_len(AsyncQueueSink_1_io_async_mem_4_len),
    .io_async_mem_4_size(AsyncQueueSink_1_io_async_mem_4_size),
    .io_async_mem_4_burst(AsyncQueueSink_1_io_async_mem_4_burst),
    .io_async_mem_4_lock(AsyncQueueSink_1_io_async_mem_4_lock),
    .io_async_mem_4_cache(AsyncQueueSink_1_io_async_mem_4_cache),
    .io_async_mem_4_prot(AsyncQueueSink_1_io_async_mem_4_prot),
    .io_async_mem_4_qos(AsyncQueueSink_1_io_async_mem_4_qos),
    .io_async_mem_5_id(AsyncQueueSink_1_io_async_mem_5_id),
    .io_async_mem_5_addr(AsyncQueueSink_1_io_async_mem_5_addr),
    .io_async_mem_5_len(AsyncQueueSink_1_io_async_mem_5_len),
    .io_async_mem_5_size(AsyncQueueSink_1_io_async_mem_5_size),
    .io_async_mem_5_burst(AsyncQueueSink_1_io_async_mem_5_burst),
    .io_async_mem_5_lock(AsyncQueueSink_1_io_async_mem_5_lock),
    .io_async_mem_5_cache(AsyncQueueSink_1_io_async_mem_5_cache),
    .io_async_mem_5_prot(AsyncQueueSink_1_io_async_mem_5_prot),
    .io_async_mem_5_qos(AsyncQueueSink_1_io_async_mem_5_qos),
    .io_async_mem_6_id(AsyncQueueSink_1_io_async_mem_6_id),
    .io_async_mem_6_addr(AsyncQueueSink_1_io_async_mem_6_addr),
    .io_async_mem_6_len(AsyncQueueSink_1_io_async_mem_6_len),
    .io_async_mem_6_size(AsyncQueueSink_1_io_async_mem_6_size),
    .io_async_mem_6_burst(AsyncQueueSink_1_io_async_mem_6_burst),
    .io_async_mem_6_lock(AsyncQueueSink_1_io_async_mem_6_lock),
    .io_async_mem_6_cache(AsyncQueueSink_1_io_async_mem_6_cache),
    .io_async_mem_6_prot(AsyncQueueSink_1_io_async_mem_6_prot),
    .io_async_mem_6_qos(AsyncQueueSink_1_io_async_mem_6_qos),
    .io_async_mem_7_id(AsyncQueueSink_1_io_async_mem_7_id),
    .io_async_mem_7_addr(AsyncQueueSink_1_io_async_mem_7_addr),
    .io_async_mem_7_len(AsyncQueueSink_1_io_async_mem_7_len),
    .io_async_mem_7_size(AsyncQueueSink_1_io_async_mem_7_size),
    .io_async_mem_7_burst(AsyncQueueSink_1_io_async_mem_7_burst),
    .io_async_mem_7_lock(AsyncQueueSink_1_io_async_mem_7_lock),
    .io_async_mem_7_cache(AsyncQueueSink_1_io_async_mem_7_cache),
    .io_async_mem_7_prot(AsyncQueueSink_1_io_async_mem_7_prot),
    .io_async_mem_7_qos(AsyncQueueSink_1_io_async_mem_7_qos),
    .io_async_ridx(AsyncQueueSink_1_io_async_ridx),
    .io_async_widx(AsyncQueueSink_1_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_1_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_1_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_1_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_1_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink_5 AsyncQueueSink_2 ( // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305085.4]
    .clock(AsyncQueueSink_2_clock),
    .reset(AsyncQueueSink_2_reset),
    .io_deq_ready(AsyncQueueSink_2_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_2_io_deq_valid),
    .io_deq_bits_data(AsyncQueueSink_2_io_deq_bits_data),
    .io_deq_bits_strb(AsyncQueueSink_2_io_deq_bits_strb),
    .io_deq_bits_last(AsyncQueueSink_2_io_deq_bits_last),
    .io_async_mem_0_data(AsyncQueueSink_2_io_async_mem_0_data),
    .io_async_mem_0_strb(AsyncQueueSink_2_io_async_mem_0_strb),
    .io_async_mem_0_last(AsyncQueueSink_2_io_async_mem_0_last),
    .io_async_mem_1_data(AsyncQueueSink_2_io_async_mem_1_data),
    .io_async_mem_1_strb(AsyncQueueSink_2_io_async_mem_1_strb),
    .io_async_mem_1_last(AsyncQueueSink_2_io_async_mem_1_last),
    .io_async_mem_2_data(AsyncQueueSink_2_io_async_mem_2_data),
    .io_async_mem_2_strb(AsyncQueueSink_2_io_async_mem_2_strb),
    .io_async_mem_2_last(AsyncQueueSink_2_io_async_mem_2_last),
    .io_async_mem_3_data(AsyncQueueSink_2_io_async_mem_3_data),
    .io_async_mem_3_strb(AsyncQueueSink_2_io_async_mem_3_strb),
    .io_async_mem_3_last(AsyncQueueSink_2_io_async_mem_3_last),
    .io_async_mem_4_data(AsyncQueueSink_2_io_async_mem_4_data),
    .io_async_mem_4_strb(AsyncQueueSink_2_io_async_mem_4_strb),
    .io_async_mem_4_last(AsyncQueueSink_2_io_async_mem_4_last),
    .io_async_mem_5_data(AsyncQueueSink_2_io_async_mem_5_data),
    .io_async_mem_5_strb(AsyncQueueSink_2_io_async_mem_5_strb),
    .io_async_mem_5_last(AsyncQueueSink_2_io_async_mem_5_last),
    .io_async_mem_6_data(AsyncQueueSink_2_io_async_mem_6_data),
    .io_async_mem_6_strb(AsyncQueueSink_2_io_async_mem_6_strb),
    .io_async_mem_6_last(AsyncQueueSink_2_io_async_mem_6_last),
    .io_async_mem_7_data(AsyncQueueSink_2_io_async_mem_7_data),
    .io_async_mem_7_strb(AsyncQueueSink_2_io_async_mem_7_strb),
    .io_async_mem_7_last(AsyncQueueSink_2_io_async_mem_7_last),
    .io_async_ridx(AsyncQueueSink_2_io_async_ridx),
    .io_async_widx(AsyncQueueSink_2_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_2_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_2_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_2_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_2_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource_3 AsyncQueueSource ( // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305103.4]
    .clock(AsyncQueueSource_clock),
    .reset(AsyncQueueSource_reset),
    .io_enq_ready(AsyncQueueSource_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_io_enq_valid),
    .io_enq_bits_id(AsyncQueueSource_io_enq_bits_id),
    .io_enq_bits_data(AsyncQueueSource_io_enq_bits_data),
    .io_enq_bits_resp(AsyncQueueSource_io_enq_bits_resp),
    .io_enq_bits_last(AsyncQueueSource_io_enq_bits_last),
    .io_async_mem_0_id(AsyncQueueSource_io_async_mem_0_id),
    .io_async_mem_0_data(AsyncQueueSource_io_async_mem_0_data),
    .io_async_mem_0_resp(AsyncQueueSource_io_async_mem_0_resp),
    .io_async_mem_0_last(AsyncQueueSource_io_async_mem_0_last),
    .io_async_mem_1_id(AsyncQueueSource_io_async_mem_1_id),
    .io_async_mem_1_data(AsyncQueueSource_io_async_mem_1_data),
    .io_async_mem_1_resp(AsyncQueueSource_io_async_mem_1_resp),
    .io_async_mem_1_last(AsyncQueueSource_io_async_mem_1_last),
    .io_async_mem_2_id(AsyncQueueSource_io_async_mem_2_id),
    .io_async_mem_2_data(AsyncQueueSource_io_async_mem_2_data),
    .io_async_mem_2_resp(AsyncQueueSource_io_async_mem_2_resp),
    .io_async_mem_2_last(AsyncQueueSource_io_async_mem_2_last),
    .io_async_mem_3_id(AsyncQueueSource_io_async_mem_3_id),
    .io_async_mem_3_data(AsyncQueueSource_io_async_mem_3_data),
    .io_async_mem_3_resp(AsyncQueueSource_io_async_mem_3_resp),
    .io_async_mem_3_last(AsyncQueueSource_io_async_mem_3_last),
    .io_async_mem_4_id(AsyncQueueSource_io_async_mem_4_id),
    .io_async_mem_4_data(AsyncQueueSource_io_async_mem_4_data),
    .io_async_mem_4_resp(AsyncQueueSource_io_async_mem_4_resp),
    .io_async_mem_4_last(AsyncQueueSource_io_async_mem_4_last),
    .io_async_mem_5_id(AsyncQueueSource_io_async_mem_5_id),
    .io_async_mem_5_data(AsyncQueueSource_io_async_mem_5_data),
    .io_async_mem_5_resp(AsyncQueueSource_io_async_mem_5_resp),
    .io_async_mem_5_last(AsyncQueueSource_io_async_mem_5_last),
    .io_async_mem_6_id(AsyncQueueSource_io_async_mem_6_id),
    .io_async_mem_6_data(AsyncQueueSource_io_async_mem_6_data),
    .io_async_mem_6_resp(AsyncQueueSource_io_async_mem_6_resp),
    .io_async_mem_6_last(AsyncQueueSource_io_async_mem_6_last),
    .io_async_mem_7_id(AsyncQueueSource_io_async_mem_7_id),
    .io_async_mem_7_data(AsyncQueueSource_io_async_mem_7_data),
    .io_async_mem_7_resp(AsyncQueueSource_io_async_mem_7_resp),
    .io_async_mem_7_last(AsyncQueueSource_io_async_mem_7_last),
    .io_async_ridx(AsyncQueueSource_io_async_ridx),
    .io_async_widx(AsyncQueueSource_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource_4 AsyncQueueSource_1 ( // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305110.4]
    .clock(AsyncQueueSource_1_clock),
    .reset(AsyncQueueSource_1_reset),
    .io_enq_ready(AsyncQueueSource_1_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_1_io_enq_valid),
    .io_enq_bits_id(AsyncQueueSource_1_io_enq_bits_id),
    .io_enq_bits_resp(AsyncQueueSource_1_io_enq_bits_resp),
    .io_async_mem_0_id(AsyncQueueSource_1_io_async_mem_0_id),
    .io_async_mem_0_resp(AsyncQueueSource_1_io_async_mem_0_resp),
    .io_async_mem_1_id(AsyncQueueSource_1_io_async_mem_1_id),
    .io_async_mem_1_resp(AsyncQueueSource_1_io_async_mem_1_resp),
    .io_async_mem_2_id(AsyncQueueSource_1_io_async_mem_2_id),
    .io_async_mem_2_resp(AsyncQueueSource_1_io_async_mem_2_resp),
    .io_async_mem_3_id(AsyncQueueSource_1_io_async_mem_3_id),
    .io_async_mem_3_resp(AsyncQueueSource_1_io_async_mem_3_resp),
    .io_async_mem_4_id(AsyncQueueSource_1_io_async_mem_4_id),
    .io_async_mem_4_resp(AsyncQueueSource_1_io_async_mem_4_resp),
    .io_async_mem_5_id(AsyncQueueSource_1_io_async_mem_5_id),
    .io_async_mem_5_resp(AsyncQueueSource_1_io_async_mem_5_resp),
    .io_async_mem_6_id(AsyncQueueSource_1_io_async_mem_6_id),
    .io_async_mem_6_resp(AsyncQueueSource_1_io_async_mem_6_resp),
    .io_async_mem_7_id(AsyncQueueSource_1_io_async_mem_7_id),
    .io_async_mem_7_resp(AsyncQueueSource_1_io_async_mem_7_resp),
    .io_async_ridx(AsyncQueueSource_1_io_async_ridx),
    .io_async_widx(AsyncQueueSource_1_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_1_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_1_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_1_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_1_io_async_safe_sink_reset_n)
  );
  assign auto_in_aw_ridx = AsyncQueueSink_1_io_async_ridx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_aw_safe_ridx_valid = AsyncQueueSink_1_io_async_safe_ridx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_aw_safe_sink_reset_n = AsyncQueueSink_1_io_async_safe_sink_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_w_ridx = AsyncQueueSink_2_io_async_ridx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_w_safe_ridx_valid = AsyncQueueSink_2_io_async_safe_ridx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_w_safe_sink_reset_n = AsyncQueueSink_2_io_async_safe_sink_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_0_id = AsyncQueueSource_1_io_async_mem_0_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_0_resp = AsyncQueueSource_1_io_async_mem_0_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_1_id = AsyncQueueSource_1_io_async_mem_1_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_1_resp = AsyncQueueSource_1_io_async_mem_1_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_2_id = AsyncQueueSource_1_io_async_mem_2_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_2_resp = AsyncQueueSource_1_io_async_mem_2_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_3_id = AsyncQueueSource_1_io_async_mem_3_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_3_resp = AsyncQueueSource_1_io_async_mem_3_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_4_id = AsyncQueueSource_1_io_async_mem_4_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_4_resp = AsyncQueueSource_1_io_async_mem_4_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_5_id = AsyncQueueSource_1_io_async_mem_5_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_5_resp = AsyncQueueSource_1_io_async_mem_5_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_6_id = AsyncQueueSource_1_io_async_mem_6_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_6_resp = AsyncQueueSource_1_io_async_mem_6_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_7_id = AsyncQueueSource_1_io_async_mem_7_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_mem_7_resp = AsyncQueueSource_1_io_async_mem_7_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_widx = AsyncQueueSource_1_io_async_widx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_safe_widx_valid = AsyncQueueSource_1_io_async_safe_widx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_b_safe_source_reset_n = AsyncQueueSource_1_io_async_safe_source_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_ar_ridx = AsyncQueueSink_io_async_ridx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_ar_safe_ridx_valid = AsyncQueueSink_io_async_safe_ridx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_ar_safe_sink_reset_n = AsyncQueueSink_io_async_safe_sink_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_0_id = AsyncQueueSource_io_async_mem_0_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_0_data = AsyncQueueSource_io_async_mem_0_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_0_resp = AsyncQueueSource_io_async_mem_0_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_0_last = AsyncQueueSource_io_async_mem_0_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_1_id = AsyncQueueSource_io_async_mem_1_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_1_data = AsyncQueueSource_io_async_mem_1_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_1_resp = AsyncQueueSource_io_async_mem_1_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_1_last = AsyncQueueSource_io_async_mem_1_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_2_id = AsyncQueueSource_io_async_mem_2_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_2_data = AsyncQueueSource_io_async_mem_2_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_2_resp = AsyncQueueSource_io_async_mem_2_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_2_last = AsyncQueueSource_io_async_mem_2_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_3_id = AsyncQueueSource_io_async_mem_3_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_3_data = AsyncQueueSource_io_async_mem_3_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_3_resp = AsyncQueueSource_io_async_mem_3_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_3_last = AsyncQueueSource_io_async_mem_3_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_4_id = AsyncQueueSource_io_async_mem_4_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_4_data = AsyncQueueSource_io_async_mem_4_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_4_resp = AsyncQueueSource_io_async_mem_4_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_4_last = AsyncQueueSource_io_async_mem_4_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_5_id = AsyncQueueSource_io_async_mem_5_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_5_data = AsyncQueueSource_io_async_mem_5_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_5_resp = AsyncQueueSource_io_async_mem_5_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_5_last = AsyncQueueSource_io_async_mem_5_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_6_id = AsyncQueueSource_io_async_mem_6_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_6_data = AsyncQueueSource_io_async_mem_6_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_6_resp = AsyncQueueSource_io_async_mem_6_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_6_last = AsyncQueueSource_io_async_mem_6_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_7_id = AsyncQueueSource_io_async_mem_7_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_7_data = AsyncQueueSource_io_async_mem_7_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_7_resp = AsyncQueueSource_io_async_mem_7_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_mem_7_last = AsyncQueueSource_io_async_mem_7_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_widx = AsyncQueueSource_io_async_widx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_safe_widx_valid = AsyncQueueSource_io_async_safe_widx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_in_r_safe_source_reset_n = AsyncQueueSource_io_async_safe_source_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305048.4]
  assign auto_out_aw_valid = AsyncQueueSink_1_io_deq_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_aw_bits_id = AsyncQueueSink_1_io_deq_bits_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_aw_bits_addr = AsyncQueueSink_1_io_deq_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_aw_bits_len = AsyncQueueSink_1_io_deq_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_aw_bits_size = AsyncQueueSink_1_io_deq_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_aw_bits_burst = AsyncQueueSink_1_io_deq_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_aw_bits_lock = AsyncQueueSink_1_io_deq_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_aw_bits_prot = AsyncQueueSink_1_io_deq_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_aw_bits_qos = AsyncQueueSink_1_io_deq_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_w_valid = AsyncQueueSink_2_io_deq_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_w_bits_data = AsyncQueueSink_2_io_deq_bits_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_w_bits_strb = AsyncQueueSink_2_io_deq_bits_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_w_bits_last = AsyncQueueSink_2_io_deq_bits_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_b_ready = AsyncQueueSource_1_io_enq_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_valid = AsyncQueueSink_io_deq_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_bits_id = AsyncQueueSink_io_deq_bits_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_bits_addr = AsyncQueueSink_io_deq_bits_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_bits_len = AsyncQueueSink_io_deq_bits_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_bits_size = AsyncQueueSink_io_deq_bits_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_bits_burst = AsyncQueueSink_io_deq_bits_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_bits_lock = AsyncQueueSink_io_deq_bits_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_bits_prot = AsyncQueueSink_io_deq_bits_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_ar_bits_qos = AsyncQueueSink_io_deq_bits_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign auto_out_r_ready = AsyncQueueSource_io_enq_ready; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305047.4]
  assign AsyncQueueSink_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305050.4]
  assign AsyncQueueSink_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305051.4]
  assign AsyncQueueSink_io_deq_ready = auto_out_ar_ready; // @[AsyncCrossing.scala 38:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305066.4]
  assign AsyncQueueSink_io_async_mem_0_id = auto_in_ar_mem_0_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_0_addr = auto_in_ar_mem_0_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_0_len = auto_in_ar_mem_0_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_0_size = auto_in_ar_mem_0_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_0_burst = auto_in_ar_mem_0_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_0_lock = auto_in_ar_mem_0_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_0_cache = auto_in_ar_mem_0_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_0_prot = auto_in_ar_mem_0_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_0_qos = auto_in_ar_mem_0_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305058.4]
  assign AsyncQueueSink_io_async_mem_1_id = auto_in_ar_mem_1_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_1_addr = auto_in_ar_mem_1_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_1_len = auto_in_ar_mem_1_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_1_size = auto_in_ar_mem_1_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_1_burst = auto_in_ar_mem_1_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_1_lock = auto_in_ar_mem_1_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_1_cache = auto_in_ar_mem_1_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_1_prot = auto_in_ar_mem_1_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_1_qos = auto_in_ar_mem_1_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305059.4]
  assign AsyncQueueSink_io_async_mem_2_id = auto_in_ar_mem_2_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_2_addr = auto_in_ar_mem_2_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_2_len = auto_in_ar_mem_2_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_2_size = auto_in_ar_mem_2_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_2_burst = auto_in_ar_mem_2_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_2_lock = auto_in_ar_mem_2_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_2_cache = auto_in_ar_mem_2_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_2_prot = auto_in_ar_mem_2_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_2_qos = auto_in_ar_mem_2_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305060.4]
  assign AsyncQueueSink_io_async_mem_3_id = auto_in_ar_mem_3_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_3_addr = auto_in_ar_mem_3_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_3_len = auto_in_ar_mem_3_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_3_size = auto_in_ar_mem_3_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_3_burst = auto_in_ar_mem_3_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_3_lock = auto_in_ar_mem_3_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_3_cache = auto_in_ar_mem_3_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_3_prot = auto_in_ar_mem_3_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_3_qos = auto_in_ar_mem_3_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305061.4]
  assign AsyncQueueSink_io_async_mem_4_id = auto_in_ar_mem_4_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_4_addr = auto_in_ar_mem_4_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_4_len = auto_in_ar_mem_4_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_4_size = auto_in_ar_mem_4_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_4_burst = auto_in_ar_mem_4_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_4_lock = auto_in_ar_mem_4_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_4_cache = auto_in_ar_mem_4_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_4_prot = auto_in_ar_mem_4_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_4_qos = auto_in_ar_mem_4_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305062.4]
  assign AsyncQueueSink_io_async_mem_5_id = auto_in_ar_mem_5_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_5_addr = auto_in_ar_mem_5_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_5_len = auto_in_ar_mem_5_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_5_size = auto_in_ar_mem_5_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_5_burst = auto_in_ar_mem_5_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_5_lock = auto_in_ar_mem_5_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_5_cache = auto_in_ar_mem_5_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_5_prot = auto_in_ar_mem_5_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_5_qos = auto_in_ar_mem_5_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305063.4]
  assign AsyncQueueSink_io_async_mem_6_id = auto_in_ar_mem_6_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_6_addr = auto_in_ar_mem_6_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_6_len = auto_in_ar_mem_6_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_6_size = auto_in_ar_mem_6_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_6_burst = auto_in_ar_mem_6_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_6_lock = auto_in_ar_mem_6_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_6_cache = auto_in_ar_mem_6_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_6_prot = auto_in_ar_mem_6_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_6_qos = auto_in_ar_mem_6_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305064.4]
  assign AsyncQueueSink_io_async_mem_7_id = auto_in_ar_mem_7_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_mem_7_addr = auto_in_ar_mem_7_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_mem_7_len = auto_in_ar_mem_7_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_mem_7_size = auto_in_ar_mem_7_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_mem_7_burst = auto_in_ar_mem_7_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_mem_7_lock = auto_in_ar_mem_7_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_mem_7_cache = auto_in_ar_mem_7_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_mem_7_prot = auto_in_ar_mem_7_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_mem_7_qos = auto_in_ar_mem_7_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305065.4]
  assign AsyncQueueSink_io_async_widx = auto_in_ar_widx; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305056.4]
  assign AsyncQueueSink_io_async_safe_widx_valid = auto_in_ar_safe_widx_valid; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305054.4]
  assign AsyncQueueSink_io_async_safe_source_reset_n = auto_in_ar_safe_source_reset_n; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305053.4]
  assign AsyncQueueSink_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305068.4]
  assign AsyncQueueSink_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305069.4]
  assign AsyncQueueSink_1_io_deq_ready = auto_out_aw_ready; // @[AsyncCrossing.scala 39:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305084.4]
  assign AsyncQueueSink_1_io_async_mem_0_id = auto_in_aw_mem_0_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_0_addr = auto_in_aw_mem_0_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_0_len = auto_in_aw_mem_0_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_0_size = auto_in_aw_mem_0_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_0_burst = auto_in_aw_mem_0_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_0_lock = auto_in_aw_mem_0_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_0_cache = auto_in_aw_mem_0_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_0_prot = auto_in_aw_mem_0_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_0_qos = auto_in_aw_mem_0_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305076.4]
  assign AsyncQueueSink_1_io_async_mem_1_id = auto_in_aw_mem_1_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_1_addr = auto_in_aw_mem_1_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_1_len = auto_in_aw_mem_1_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_1_size = auto_in_aw_mem_1_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_1_burst = auto_in_aw_mem_1_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_1_lock = auto_in_aw_mem_1_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_1_cache = auto_in_aw_mem_1_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_1_prot = auto_in_aw_mem_1_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_1_qos = auto_in_aw_mem_1_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305077.4]
  assign AsyncQueueSink_1_io_async_mem_2_id = auto_in_aw_mem_2_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_2_addr = auto_in_aw_mem_2_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_2_len = auto_in_aw_mem_2_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_2_size = auto_in_aw_mem_2_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_2_burst = auto_in_aw_mem_2_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_2_lock = auto_in_aw_mem_2_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_2_cache = auto_in_aw_mem_2_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_2_prot = auto_in_aw_mem_2_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_2_qos = auto_in_aw_mem_2_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305078.4]
  assign AsyncQueueSink_1_io_async_mem_3_id = auto_in_aw_mem_3_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_3_addr = auto_in_aw_mem_3_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_3_len = auto_in_aw_mem_3_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_3_size = auto_in_aw_mem_3_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_3_burst = auto_in_aw_mem_3_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_3_lock = auto_in_aw_mem_3_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_3_cache = auto_in_aw_mem_3_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_3_prot = auto_in_aw_mem_3_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_3_qos = auto_in_aw_mem_3_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305079.4]
  assign AsyncQueueSink_1_io_async_mem_4_id = auto_in_aw_mem_4_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_4_addr = auto_in_aw_mem_4_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_4_len = auto_in_aw_mem_4_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_4_size = auto_in_aw_mem_4_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_4_burst = auto_in_aw_mem_4_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_4_lock = auto_in_aw_mem_4_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_4_cache = auto_in_aw_mem_4_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_4_prot = auto_in_aw_mem_4_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_4_qos = auto_in_aw_mem_4_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305080.4]
  assign AsyncQueueSink_1_io_async_mem_5_id = auto_in_aw_mem_5_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_5_addr = auto_in_aw_mem_5_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_5_len = auto_in_aw_mem_5_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_5_size = auto_in_aw_mem_5_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_5_burst = auto_in_aw_mem_5_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_5_lock = auto_in_aw_mem_5_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_5_cache = auto_in_aw_mem_5_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_5_prot = auto_in_aw_mem_5_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_5_qos = auto_in_aw_mem_5_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305081.4]
  assign AsyncQueueSink_1_io_async_mem_6_id = auto_in_aw_mem_6_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_6_addr = auto_in_aw_mem_6_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_6_len = auto_in_aw_mem_6_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_6_size = auto_in_aw_mem_6_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_6_burst = auto_in_aw_mem_6_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_6_lock = auto_in_aw_mem_6_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_6_cache = auto_in_aw_mem_6_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_6_prot = auto_in_aw_mem_6_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_6_qos = auto_in_aw_mem_6_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305082.4]
  assign AsyncQueueSink_1_io_async_mem_7_id = auto_in_aw_mem_7_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_mem_7_addr = auto_in_aw_mem_7_addr; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_mem_7_len = auto_in_aw_mem_7_len; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_mem_7_size = auto_in_aw_mem_7_size; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_mem_7_burst = auto_in_aw_mem_7_burst; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_mem_7_lock = auto_in_aw_mem_7_lock; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_mem_7_cache = auto_in_aw_mem_7_cache; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_mem_7_prot = auto_in_aw_mem_7_prot; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_mem_7_qos = auto_in_aw_mem_7_qos; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305083.4]
  assign AsyncQueueSink_1_io_async_widx = auto_in_aw_widx; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305074.4]
  assign AsyncQueueSink_1_io_async_safe_widx_valid = auto_in_aw_safe_widx_valid; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305072.4]
  assign AsyncQueueSink_1_io_async_safe_source_reset_n = auto_in_aw_safe_source_reset_n; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305071.4]
  assign AsyncQueueSink_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305086.4]
  assign AsyncQueueSink_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305087.4]
  assign AsyncQueueSink_2_io_deq_ready = auto_out_w_ready; // @[AsyncCrossing.scala 40:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305102.4]
  assign AsyncQueueSink_2_io_async_mem_0_data = auto_in_w_mem_0_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305094.4]
  assign AsyncQueueSink_2_io_async_mem_0_strb = auto_in_w_mem_0_strb; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305094.4]
  assign AsyncQueueSink_2_io_async_mem_0_last = auto_in_w_mem_0_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305094.4]
  assign AsyncQueueSink_2_io_async_mem_1_data = auto_in_w_mem_1_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305095.4]
  assign AsyncQueueSink_2_io_async_mem_1_strb = auto_in_w_mem_1_strb; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305095.4]
  assign AsyncQueueSink_2_io_async_mem_1_last = auto_in_w_mem_1_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305095.4]
  assign AsyncQueueSink_2_io_async_mem_2_data = auto_in_w_mem_2_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305096.4]
  assign AsyncQueueSink_2_io_async_mem_2_strb = auto_in_w_mem_2_strb; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305096.4]
  assign AsyncQueueSink_2_io_async_mem_2_last = auto_in_w_mem_2_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305096.4]
  assign AsyncQueueSink_2_io_async_mem_3_data = auto_in_w_mem_3_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305097.4]
  assign AsyncQueueSink_2_io_async_mem_3_strb = auto_in_w_mem_3_strb; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305097.4]
  assign AsyncQueueSink_2_io_async_mem_3_last = auto_in_w_mem_3_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305097.4]
  assign AsyncQueueSink_2_io_async_mem_4_data = auto_in_w_mem_4_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305098.4]
  assign AsyncQueueSink_2_io_async_mem_4_strb = auto_in_w_mem_4_strb; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305098.4]
  assign AsyncQueueSink_2_io_async_mem_4_last = auto_in_w_mem_4_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305098.4]
  assign AsyncQueueSink_2_io_async_mem_5_data = auto_in_w_mem_5_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305099.4]
  assign AsyncQueueSink_2_io_async_mem_5_strb = auto_in_w_mem_5_strb; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305099.4]
  assign AsyncQueueSink_2_io_async_mem_5_last = auto_in_w_mem_5_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305099.4]
  assign AsyncQueueSink_2_io_async_mem_6_data = auto_in_w_mem_6_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305100.4]
  assign AsyncQueueSink_2_io_async_mem_6_strb = auto_in_w_mem_6_strb; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305100.4]
  assign AsyncQueueSink_2_io_async_mem_6_last = auto_in_w_mem_6_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305100.4]
  assign AsyncQueueSink_2_io_async_mem_7_data = auto_in_w_mem_7_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305101.4]
  assign AsyncQueueSink_2_io_async_mem_7_strb = auto_in_w_mem_7_strb; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305101.4]
  assign AsyncQueueSink_2_io_async_mem_7_last = auto_in_w_mem_7_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305101.4]
  assign AsyncQueueSink_2_io_async_widx = auto_in_w_widx; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305092.4]
  assign AsyncQueueSink_2_io_async_safe_widx_valid = auto_in_w_safe_widx_valid; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305090.4]
  assign AsyncQueueSink_2_io_async_safe_source_reset_n = auto_in_w_safe_source_reset_n; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305089.4]
  assign AsyncQueueSource_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305104.4]
  assign AsyncQueueSource_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305105.4]
  assign AsyncQueueSource_io_enq_valid = auto_out_r_valid; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305107.4]
  assign AsyncQueueSource_io_enq_bits_id = auto_out_r_bits_id; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305106.4]
  assign AsyncQueueSource_io_enq_bits_data = auto_out_r_bits_data; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305106.4]
  assign AsyncQueueSource_io_enq_bits_resp = auto_out_r_bits_resp; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305106.4]
  assign AsyncQueueSource_io_enq_bits_last = auto_out_r_bits_last; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305106.4]
  assign AsyncQueueSource_io_async_ridx = auto_in_r_ridx; // @[AsyncCrossing.scala 41:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305109.4]
  assign AsyncQueueSource_io_async_safe_ridx_valid = auto_in_r_safe_ridx_valid; // @[AsyncCrossing.scala 41:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305109.4]
  assign AsyncQueueSource_io_async_safe_sink_reset_n = auto_in_r_safe_sink_reset_n; // @[AsyncCrossing.scala 41:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305109.4]
  assign AsyncQueueSource_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305111.4]
  assign AsyncQueueSource_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305112.4]
  assign AsyncQueueSource_1_io_enq_valid = auto_out_b_valid; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305114.4]
  assign AsyncQueueSource_1_io_enq_bits_id = auto_out_b_bits_id; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305113.4]
  assign AsyncQueueSource_1_io_enq_bits_resp = auto_out_b_bits_resp; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305113.4]
  assign AsyncQueueSource_1_io_async_ridx = auto_in_b_ridx; // @[AsyncCrossing.scala 42:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305116.4]
  assign AsyncQueueSource_1_io_async_safe_ridx_valid = auto_in_b_safe_ridx_valid; // @[AsyncCrossing.scala 42:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305116.4]
  assign AsyncQueueSource_1_io_async_safe_sink_reset_n = auto_in_b_safe_sink_reset_n; // @[AsyncCrossing.scala 42:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305116.4]
endmodule
module XilinxVC707MIGIsland( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305189.2]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_aw_mem_0_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_aw_mem_0_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_0_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_aw_mem_0_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_mem_0_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_0_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_0_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_0_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_aw_mem_1_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_aw_mem_1_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_1_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_aw_mem_1_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_mem_1_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_1_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_1_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_1_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_aw_mem_2_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_aw_mem_2_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_2_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_aw_mem_2_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_mem_2_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_2_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_2_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_2_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_aw_mem_3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_aw_mem_3_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_3_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_aw_mem_3_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_mem_3_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_3_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_3_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_3_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_aw_mem_4_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_aw_mem_4_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_4_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_aw_mem_4_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_mem_4_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_4_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_4_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_4_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_aw_mem_5_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_aw_mem_5_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_5_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_aw_mem_5_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_mem_5_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_5_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_5_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_5_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_aw_mem_6_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_aw_mem_6_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_6_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_aw_mem_6_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_mem_6_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_6_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_6_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_6_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_aw_mem_7_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_aw_mem_7_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_7_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_aw_mem_7_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_mem_7_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_7_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_aw_mem_7_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_mem_7_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_aw_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_aw_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_aw_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_aw_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_aw_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [63:0] auto_axi4in_xing_in_w_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_w_mem_0_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [63:0] auto_axi4in_xing_in_w_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_w_mem_1_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [63:0] auto_axi4in_xing_in_w_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_w_mem_2_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [63:0] auto_axi4in_xing_in_w_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_w_mem_3_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [63:0] auto_axi4in_xing_in_w_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_w_mem_4_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [63:0] auto_axi4in_xing_in_w_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_w_mem_5_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [63:0] auto_axi4in_xing_in_w_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_w_mem_6_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [63:0] auto_axi4in_xing_in_w_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_w_mem_7_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_w_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_w_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_w_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_w_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_w_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_b_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_b_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_b_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_b_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_b_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_b_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_b_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_b_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_b_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_b_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_b_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_b_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_b_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_b_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_ar_mem_0_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_ar_mem_0_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_0_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_ar_mem_0_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_mem_0_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_0_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_0_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_0_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_ar_mem_1_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_ar_mem_1_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_1_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_ar_mem_1_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_mem_1_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_1_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_1_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_1_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_ar_mem_2_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_ar_mem_2_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_2_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_ar_mem_2_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_mem_2_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_2_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_2_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_2_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_ar_mem_3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_ar_mem_3_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_3_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_ar_mem_3_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_mem_3_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_3_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_3_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_3_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_ar_mem_4_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_ar_mem_4_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_4_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_ar_mem_4_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_mem_4_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_4_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_4_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_4_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_ar_mem_5_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_ar_mem_5_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_5_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_ar_mem_5_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_mem_5_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_5_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_5_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_5_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_ar_mem_6_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_ar_mem_6_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_6_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_ar_mem_6_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_mem_6_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_6_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_6_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_6_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [31:0] auto_axi4in_xing_in_ar_mem_7_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [7:0]  auto_axi4in_xing_in_ar_mem_7_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_7_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [1:0]  auto_axi4in_xing_in_ar_mem_7_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_mem_7_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_7_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [2:0]  auto_axi4in_xing_in_ar_mem_7_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_mem_7_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_ar_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_ar_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_ar_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_ar_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_ar_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [63:0] auto_axi4in_xing_in_r_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_r_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [63:0] auto_axi4in_xing_in_r_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_r_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [63:0] auto_axi4in_xing_in_r_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_r_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [63:0] auto_axi4in_xing_in_r_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_r_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [63:0] auto_axi4in_xing_in_r_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_r_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [63:0] auto_axi4in_xing_in_r_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_r_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [63:0] auto_axi4in_xing_in_r_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_r_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [63:0] auto_axi4in_xing_in_r_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [1:0]  auto_axi4in_xing_in_r_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input  [3:0]  auto_axi4in_xing_in_r_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [3:0]  auto_axi4in_xing_in_r_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_r_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output        auto_axi4in_xing_in_r_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  input         auto_axi4in_xing_in_r_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305190.4]
  output [13:0] io_port_ddr3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output [2:0]  io_port_ddr3_ba, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_ras_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_cas_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_we_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_ck_p, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_ck_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_cke, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_cs_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output [7:0]  io_port_ddr3_dm, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ddr3_odt, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  inout  [63:0] io_port_ddr3_dq, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  inout  [7:0]  io_port_ddr3_dqs_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  inout  [7:0]  io_port_ddr3_dqs_p, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  input         io_port_sys_clk_i, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ui_clk, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_ui_clk_sync_rst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  output        io_port_mmcm_locked, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  input         io_port_aresetn, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
  input         io_port_sys_rst // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305191.4]
);
  wire  axi4asink_clock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_reset; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_0_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_aw_mem_0_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_aw_mem_0_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_0_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_aw_mem_0_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_mem_0_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_0_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_0_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_0_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_1_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_aw_mem_1_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_aw_mem_1_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_1_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_aw_mem_1_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_mem_1_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_1_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_1_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_1_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_2_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_aw_mem_2_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_aw_mem_2_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_2_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_aw_mem_2_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_mem_2_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_2_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_2_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_2_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_3_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_aw_mem_3_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_aw_mem_3_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_3_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_aw_mem_3_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_mem_3_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_3_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_3_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_3_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_4_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_aw_mem_4_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_aw_mem_4_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_4_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_aw_mem_4_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_mem_4_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_4_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_4_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_4_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_5_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_aw_mem_5_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_aw_mem_5_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_5_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_aw_mem_5_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_mem_5_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_5_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_5_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_5_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_6_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_aw_mem_6_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_aw_mem_6_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_6_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_aw_mem_6_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_mem_6_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_6_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_6_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_6_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_7_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_aw_mem_7_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_aw_mem_7_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_7_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_aw_mem_7_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_mem_7_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_7_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_aw_mem_7_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_mem_7_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_ridx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_aw_widx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_safe_ridx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_safe_widx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_safe_source_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_aw_safe_sink_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_w_mem_0_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_w_mem_0_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_mem_0_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_w_mem_1_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_w_mem_1_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_mem_1_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_w_mem_2_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_w_mem_2_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_mem_2_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_w_mem_3_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_w_mem_3_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_mem_3_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_w_mem_4_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_w_mem_4_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_mem_4_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_w_mem_5_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_w_mem_5_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_mem_5_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_w_mem_6_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_w_mem_6_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_mem_6_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_w_mem_7_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_w_mem_7_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_mem_7_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_w_ridx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_w_widx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_safe_ridx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_safe_widx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_safe_source_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_w_safe_sink_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_mem_0_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_b_mem_0_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_mem_1_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_b_mem_1_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_mem_2_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_b_mem_2_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_mem_3_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_b_mem_3_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_mem_4_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_b_mem_4_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_mem_5_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_b_mem_5_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_mem_6_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_b_mem_6_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_mem_7_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_b_mem_7_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_ridx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_b_widx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_b_safe_ridx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_b_safe_widx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_b_safe_source_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_b_safe_sink_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_0_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_ar_mem_0_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_ar_mem_0_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_0_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_ar_mem_0_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_mem_0_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_0_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_0_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_0_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_1_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_ar_mem_1_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_ar_mem_1_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_1_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_ar_mem_1_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_mem_1_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_1_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_1_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_1_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_2_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_ar_mem_2_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_ar_mem_2_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_2_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_ar_mem_2_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_mem_2_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_2_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_2_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_2_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_3_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_ar_mem_3_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_ar_mem_3_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_3_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_ar_mem_3_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_mem_3_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_3_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_3_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_3_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_4_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_ar_mem_4_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_ar_mem_4_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_4_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_ar_mem_4_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_mem_4_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_4_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_4_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_4_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_5_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_ar_mem_5_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_ar_mem_5_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_5_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_ar_mem_5_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_mem_5_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_5_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_5_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_5_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_6_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_ar_mem_6_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_ar_mem_6_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_6_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_ar_mem_6_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_mem_6_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_6_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_6_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_6_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_7_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_in_ar_mem_7_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_in_ar_mem_7_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_7_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_ar_mem_7_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_mem_7_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_7_cache; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_in_ar_mem_7_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_mem_7_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_ridx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_ar_widx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_safe_ridx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_safe_widx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_safe_source_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_ar_safe_sink_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_mem_0_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_r_mem_0_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_r_mem_0_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_mem_0_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_mem_1_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_r_mem_1_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_r_mem_1_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_mem_1_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_mem_2_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_r_mem_2_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_r_mem_2_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_mem_2_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_mem_3_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_r_mem_3_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_r_mem_3_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_mem_3_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_mem_4_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_r_mem_4_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_r_mem_4_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_mem_4_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_mem_5_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_r_mem_5_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_r_mem_5_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_mem_5_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_mem_6_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_r_mem_6_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_r_mem_6_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_mem_6_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_mem_7_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_in_r_mem_7_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_in_r_mem_7_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_mem_7_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_ridx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_in_r_widx; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_safe_ridx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_safe_widx_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_safe_source_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_in_r_safe_sink_reset_n; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_aw_ready; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_aw_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_out_aw_bits_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_out_aw_bits_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_out_aw_bits_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_out_aw_bits_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_out_aw_bits_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_aw_bits_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_out_aw_bits_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_out_aw_bits_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_w_ready; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_w_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_out_w_bits_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_out_w_bits_strb; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_w_bits_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_b_ready; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_b_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_out_b_bits_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_out_b_bits_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_ar_ready; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_ar_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_out_ar_bits_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [31:0] axi4asink_auto_out_ar_bits_addr; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [7:0] axi4asink_auto_out_ar_bits_len; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_out_ar_bits_size; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_out_ar_bits_burst; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_ar_bits_lock; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [2:0] axi4asink_auto_out_ar_bits_prot; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_out_ar_bits_qos; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_r_ready; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_r_valid; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [3:0] axi4asink_auto_out_r_bits_id; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [63:0] axi4asink_auto_out_r_bits_data; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [1:0] axi4asink_auto_out_r_bits_resp; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire  axi4asink_auto_out_r_bits_last; // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
  wire [11:0] blackbox_device_temp; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_rvalid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_rlast; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [1:0] blackbox_s_axi_rresp; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [63:0] blackbox_s_axi_rdata; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [3:0] blackbox_s_axi_rid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_rready; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_arready; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_arvalid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [3:0] blackbox_s_axi_arqos; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [2:0] blackbox_s_axi_arprot; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [3:0] blackbox_s_axi_arcache; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_arlock; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [1:0] blackbox_s_axi_arburst; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [2:0] blackbox_s_axi_arsize; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [7:0] blackbox_s_axi_arlen; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [29:0] blackbox_s_axi_araddr; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [3:0] blackbox_s_axi_arid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_bvalid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [1:0] blackbox_s_axi_bresp; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [3:0] blackbox_s_axi_bid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_bready; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_wready; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_wvalid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_wlast; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [7:0] blackbox_s_axi_wstrb; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [63:0] blackbox_s_axi_wdata; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_awready; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_awvalid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [3:0] blackbox_s_axi_awqos; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [2:0] blackbox_s_axi_awprot; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [3:0] blackbox_s_axi_awcache; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_s_axi_awlock; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [1:0] blackbox_s_axi_awburst; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [2:0] blackbox_s_axi_awsize; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [7:0] blackbox_s_axi_awlen; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [29:0] blackbox_s_axi_awaddr; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [3:0] blackbox_s_axi_awid; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_app_zq_ack; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_app_ref_ack; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_app_sr_active; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_app_zq_req; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_app_ref_req; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_app_sr_req; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_sys_rst; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_init_calib_complete; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_aresetn; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_mmcm_locked; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ui_clk_sync_rst; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ui_clk; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_sys_clk_i; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_odt; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [7:0] blackbox_ddr3_dm; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_cs_n; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_cke; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_ck_n; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_ck_p; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_reset_n; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_we_n; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_cas_n; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire  blackbox_ddr3_ras_n; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [2:0] blackbox_ddr3_ba; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [13:0] blackbox_ddr3_addr; // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
  wire [31:0] axi_async_aw_bits_addr; // @[Nodes.scala 333:76:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305208.4 LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  wire [32:0] _T_1172; // @[XilinxVC707MIG.scala 92:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305310.4]
  wire [32:0] _T_1173; // @[XilinxVC707MIG.scala 92:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305311.4]
  wire [31:0] awaddr; // @[XilinxVC707MIG.scala 92:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305312.4]
  wire [31:0] axi_async_ar_bits_addr; // @[Nodes.scala 333:76:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305208.4 LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  wire [32:0] _T_1174; // @[XilinxVC707MIG.scala 93:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305313.4]
  wire [32:0] _T_1175; // @[XilinxVC707MIG.scala 93:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305314.4]
  wire [31:0] araddr; // @[XilinxVC707MIG.scala 93:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305315.4]
  AXI4AsyncCrossingSink axi4asink ( // @[AsyncCrossing.scala 60:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305202.4]
    .clock(axi4asink_clock),
    .reset(axi4asink_reset),
    .auto_in_aw_mem_0_id(axi4asink_auto_in_aw_mem_0_id),
    .auto_in_aw_mem_0_addr(axi4asink_auto_in_aw_mem_0_addr),
    .auto_in_aw_mem_0_len(axi4asink_auto_in_aw_mem_0_len),
    .auto_in_aw_mem_0_size(axi4asink_auto_in_aw_mem_0_size),
    .auto_in_aw_mem_0_burst(axi4asink_auto_in_aw_mem_0_burst),
    .auto_in_aw_mem_0_lock(axi4asink_auto_in_aw_mem_0_lock),
    .auto_in_aw_mem_0_cache(axi4asink_auto_in_aw_mem_0_cache),
    .auto_in_aw_mem_0_prot(axi4asink_auto_in_aw_mem_0_prot),
    .auto_in_aw_mem_0_qos(axi4asink_auto_in_aw_mem_0_qos),
    .auto_in_aw_mem_1_id(axi4asink_auto_in_aw_mem_1_id),
    .auto_in_aw_mem_1_addr(axi4asink_auto_in_aw_mem_1_addr),
    .auto_in_aw_mem_1_len(axi4asink_auto_in_aw_mem_1_len),
    .auto_in_aw_mem_1_size(axi4asink_auto_in_aw_mem_1_size),
    .auto_in_aw_mem_1_burst(axi4asink_auto_in_aw_mem_1_burst),
    .auto_in_aw_mem_1_lock(axi4asink_auto_in_aw_mem_1_lock),
    .auto_in_aw_mem_1_cache(axi4asink_auto_in_aw_mem_1_cache),
    .auto_in_aw_mem_1_prot(axi4asink_auto_in_aw_mem_1_prot),
    .auto_in_aw_mem_1_qos(axi4asink_auto_in_aw_mem_1_qos),
    .auto_in_aw_mem_2_id(axi4asink_auto_in_aw_mem_2_id),
    .auto_in_aw_mem_2_addr(axi4asink_auto_in_aw_mem_2_addr),
    .auto_in_aw_mem_2_len(axi4asink_auto_in_aw_mem_2_len),
    .auto_in_aw_mem_2_size(axi4asink_auto_in_aw_mem_2_size),
    .auto_in_aw_mem_2_burst(axi4asink_auto_in_aw_mem_2_burst),
    .auto_in_aw_mem_2_lock(axi4asink_auto_in_aw_mem_2_lock),
    .auto_in_aw_mem_2_cache(axi4asink_auto_in_aw_mem_2_cache),
    .auto_in_aw_mem_2_prot(axi4asink_auto_in_aw_mem_2_prot),
    .auto_in_aw_mem_2_qos(axi4asink_auto_in_aw_mem_2_qos),
    .auto_in_aw_mem_3_id(axi4asink_auto_in_aw_mem_3_id),
    .auto_in_aw_mem_3_addr(axi4asink_auto_in_aw_mem_3_addr),
    .auto_in_aw_mem_3_len(axi4asink_auto_in_aw_mem_3_len),
    .auto_in_aw_mem_3_size(axi4asink_auto_in_aw_mem_3_size),
    .auto_in_aw_mem_3_burst(axi4asink_auto_in_aw_mem_3_burst),
    .auto_in_aw_mem_3_lock(axi4asink_auto_in_aw_mem_3_lock),
    .auto_in_aw_mem_3_cache(axi4asink_auto_in_aw_mem_3_cache),
    .auto_in_aw_mem_3_prot(axi4asink_auto_in_aw_mem_3_prot),
    .auto_in_aw_mem_3_qos(axi4asink_auto_in_aw_mem_3_qos),
    .auto_in_aw_mem_4_id(axi4asink_auto_in_aw_mem_4_id),
    .auto_in_aw_mem_4_addr(axi4asink_auto_in_aw_mem_4_addr),
    .auto_in_aw_mem_4_len(axi4asink_auto_in_aw_mem_4_len),
    .auto_in_aw_mem_4_size(axi4asink_auto_in_aw_mem_4_size),
    .auto_in_aw_mem_4_burst(axi4asink_auto_in_aw_mem_4_burst),
    .auto_in_aw_mem_4_lock(axi4asink_auto_in_aw_mem_4_lock),
    .auto_in_aw_mem_4_cache(axi4asink_auto_in_aw_mem_4_cache),
    .auto_in_aw_mem_4_prot(axi4asink_auto_in_aw_mem_4_prot),
    .auto_in_aw_mem_4_qos(axi4asink_auto_in_aw_mem_4_qos),
    .auto_in_aw_mem_5_id(axi4asink_auto_in_aw_mem_5_id),
    .auto_in_aw_mem_5_addr(axi4asink_auto_in_aw_mem_5_addr),
    .auto_in_aw_mem_5_len(axi4asink_auto_in_aw_mem_5_len),
    .auto_in_aw_mem_5_size(axi4asink_auto_in_aw_mem_5_size),
    .auto_in_aw_mem_5_burst(axi4asink_auto_in_aw_mem_5_burst),
    .auto_in_aw_mem_5_lock(axi4asink_auto_in_aw_mem_5_lock),
    .auto_in_aw_mem_5_cache(axi4asink_auto_in_aw_mem_5_cache),
    .auto_in_aw_mem_5_prot(axi4asink_auto_in_aw_mem_5_prot),
    .auto_in_aw_mem_5_qos(axi4asink_auto_in_aw_mem_5_qos),
    .auto_in_aw_mem_6_id(axi4asink_auto_in_aw_mem_6_id),
    .auto_in_aw_mem_6_addr(axi4asink_auto_in_aw_mem_6_addr),
    .auto_in_aw_mem_6_len(axi4asink_auto_in_aw_mem_6_len),
    .auto_in_aw_mem_6_size(axi4asink_auto_in_aw_mem_6_size),
    .auto_in_aw_mem_6_burst(axi4asink_auto_in_aw_mem_6_burst),
    .auto_in_aw_mem_6_lock(axi4asink_auto_in_aw_mem_6_lock),
    .auto_in_aw_mem_6_cache(axi4asink_auto_in_aw_mem_6_cache),
    .auto_in_aw_mem_6_prot(axi4asink_auto_in_aw_mem_6_prot),
    .auto_in_aw_mem_6_qos(axi4asink_auto_in_aw_mem_6_qos),
    .auto_in_aw_mem_7_id(axi4asink_auto_in_aw_mem_7_id),
    .auto_in_aw_mem_7_addr(axi4asink_auto_in_aw_mem_7_addr),
    .auto_in_aw_mem_7_len(axi4asink_auto_in_aw_mem_7_len),
    .auto_in_aw_mem_7_size(axi4asink_auto_in_aw_mem_7_size),
    .auto_in_aw_mem_7_burst(axi4asink_auto_in_aw_mem_7_burst),
    .auto_in_aw_mem_7_lock(axi4asink_auto_in_aw_mem_7_lock),
    .auto_in_aw_mem_7_cache(axi4asink_auto_in_aw_mem_7_cache),
    .auto_in_aw_mem_7_prot(axi4asink_auto_in_aw_mem_7_prot),
    .auto_in_aw_mem_7_qos(axi4asink_auto_in_aw_mem_7_qos),
    .auto_in_aw_ridx(axi4asink_auto_in_aw_ridx),
    .auto_in_aw_widx(axi4asink_auto_in_aw_widx),
    .auto_in_aw_safe_ridx_valid(axi4asink_auto_in_aw_safe_ridx_valid),
    .auto_in_aw_safe_widx_valid(axi4asink_auto_in_aw_safe_widx_valid),
    .auto_in_aw_safe_source_reset_n(axi4asink_auto_in_aw_safe_source_reset_n),
    .auto_in_aw_safe_sink_reset_n(axi4asink_auto_in_aw_safe_sink_reset_n),
    .auto_in_w_mem_0_data(axi4asink_auto_in_w_mem_0_data),
    .auto_in_w_mem_0_strb(axi4asink_auto_in_w_mem_0_strb),
    .auto_in_w_mem_0_last(axi4asink_auto_in_w_mem_0_last),
    .auto_in_w_mem_1_data(axi4asink_auto_in_w_mem_1_data),
    .auto_in_w_mem_1_strb(axi4asink_auto_in_w_mem_1_strb),
    .auto_in_w_mem_1_last(axi4asink_auto_in_w_mem_1_last),
    .auto_in_w_mem_2_data(axi4asink_auto_in_w_mem_2_data),
    .auto_in_w_mem_2_strb(axi4asink_auto_in_w_mem_2_strb),
    .auto_in_w_mem_2_last(axi4asink_auto_in_w_mem_2_last),
    .auto_in_w_mem_3_data(axi4asink_auto_in_w_mem_3_data),
    .auto_in_w_mem_3_strb(axi4asink_auto_in_w_mem_3_strb),
    .auto_in_w_mem_3_last(axi4asink_auto_in_w_mem_3_last),
    .auto_in_w_mem_4_data(axi4asink_auto_in_w_mem_4_data),
    .auto_in_w_mem_4_strb(axi4asink_auto_in_w_mem_4_strb),
    .auto_in_w_mem_4_last(axi4asink_auto_in_w_mem_4_last),
    .auto_in_w_mem_5_data(axi4asink_auto_in_w_mem_5_data),
    .auto_in_w_mem_5_strb(axi4asink_auto_in_w_mem_5_strb),
    .auto_in_w_mem_5_last(axi4asink_auto_in_w_mem_5_last),
    .auto_in_w_mem_6_data(axi4asink_auto_in_w_mem_6_data),
    .auto_in_w_mem_6_strb(axi4asink_auto_in_w_mem_6_strb),
    .auto_in_w_mem_6_last(axi4asink_auto_in_w_mem_6_last),
    .auto_in_w_mem_7_data(axi4asink_auto_in_w_mem_7_data),
    .auto_in_w_mem_7_strb(axi4asink_auto_in_w_mem_7_strb),
    .auto_in_w_mem_7_last(axi4asink_auto_in_w_mem_7_last),
    .auto_in_w_ridx(axi4asink_auto_in_w_ridx),
    .auto_in_w_widx(axi4asink_auto_in_w_widx),
    .auto_in_w_safe_ridx_valid(axi4asink_auto_in_w_safe_ridx_valid),
    .auto_in_w_safe_widx_valid(axi4asink_auto_in_w_safe_widx_valid),
    .auto_in_w_safe_source_reset_n(axi4asink_auto_in_w_safe_source_reset_n),
    .auto_in_w_safe_sink_reset_n(axi4asink_auto_in_w_safe_sink_reset_n),
    .auto_in_b_mem_0_id(axi4asink_auto_in_b_mem_0_id),
    .auto_in_b_mem_0_resp(axi4asink_auto_in_b_mem_0_resp),
    .auto_in_b_mem_1_id(axi4asink_auto_in_b_mem_1_id),
    .auto_in_b_mem_1_resp(axi4asink_auto_in_b_mem_1_resp),
    .auto_in_b_mem_2_id(axi4asink_auto_in_b_mem_2_id),
    .auto_in_b_mem_2_resp(axi4asink_auto_in_b_mem_2_resp),
    .auto_in_b_mem_3_id(axi4asink_auto_in_b_mem_3_id),
    .auto_in_b_mem_3_resp(axi4asink_auto_in_b_mem_3_resp),
    .auto_in_b_mem_4_id(axi4asink_auto_in_b_mem_4_id),
    .auto_in_b_mem_4_resp(axi4asink_auto_in_b_mem_4_resp),
    .auto_in_b_mem_5_id(axi4asink_auto_in_b_mem_5_id),
    .auto_in_b_mem_5_resp(axi4asink_auto_in_b_mem_5_resp),
    .auto_in_b_mem_6_id(axi4asink_auto_in_b_mem_6_id),
    .auto_in_b_mem_6_resp(axi4asink_auto_in_b_mem_6_resp),
    .auto_in_b_mem_7_id(axi4asink_auto_in_b_mem_7_id),
    .auto_in_b_mem_7_resp(axi4asink_auto_in_b_mem_7_resp),
    .auto_in_b_ridx(axi4asink_auto_in_b_ridx),
    .auto_in_b_widx(axi4asink_auto_in_b_widx),
    .auto_in_b_safe_ridx_valid(axi4asink_auto_in_b_safe_ridx_valid),
    .auto_in_b_safe_widx_valid(axi4asink_auto_in_b_safe_widx_valid),
    .auto_in_b_safe_source_reset_n(axi4asink_auto_in_b_safe_source_reset_n),
    .auto_in_b_safe_sink_reset_n(axi4asink_auto_in_b_safe_sink_reset_n),
    .auto_in_ar_mem_0_id(axi4asink_auto_in_ar_mem_0_id),
    .auto_in_ar_mem_0_addr(axi4asink_auto_in_ar_mem_0_addr),
    .auto_in_ar_mem_0_len(axi4asink_auto_in_ar_mem_0_len),
    .auto_in_ar_mem_0_size(axi4asink_auto_in_ar_mem_0_size),
    .auto_in_ar_mem_0_burst(axi4asink_auto_in_ar_mem_0_burst),
    .auto_in_ar_mem_0_lock(axi4asink_auto_in_ar_mem_0_lock),
    .auto_in_ar_mem_0_cache(axi4asink_auto_in_ar_mem_0_cache),
    .auto_in_ar_mem_0_prot(axi4asink_auto_in_ar_mem_0_prot),
    .auto_in_ar_mem_0_qos(axi4asink_auto_in_ar_mem_0_qos),
    .auto_in_ar_mem_1_id(axi4asink_auto_in_ar_mem_1_id),
    .auto_in_ar_mem_1_addr(axi4asink_auto_in_ar_mem_1_addr),
    .auto_in_ar_mem_1_len(axi4asink_auto_in_ar_mem_1_len),
    .auto_in_ar_mem_1_size(axi4asink_auto_in_ar_mem_1_size),
    .auto_in_ar_mem_1_burst(axi4asink_auto_in_ar_mem_1_burst),
    .auto_in_ar_mem_1_lock(axi4asink_auto_in_ar_mem_1_lock),
    .auto_in_ar_mem_1_cache(axi4asink_auto_in_ar_mem_1_cache),
    .auto_in_ar_mem_1_prot(axi4asink_auto_in_ar_mem_1_prot),
    .auto_in_ar_mem_1_qos(axi4asink_auto_in_ar_mem_1_qos),
    .auto_in_ar_mem_2_id(axi4asink_auto_in_ar_mem_2_id),
    .auto_in_ar_mem_2_addr(axi4asink_auto_in_ar_mem_2_addr),
    .auto_in_ar_mem_2_len(axi4asink_auto_in_ar_mem_2_len),
    .auto_in_ar_mem_2_size(axi4asink_auto_in_ar_mem_2_size),
    .auto_in_ar_mem_2_burst(axi4asink_auto_in_ar_mem_2_burst),
    .auto_in_ar_mem_2_lock(axi4asink_auto_in_ar_mem_2_lock),
    .auto_in_ar_mem_2_cache(axi4asink_auto_in_ar_mem_2_cache),
    .auto_in_ar_mem_2_prot(axi4asink_auto_in_ar_mem_2_prot),
    .auto_in_ar_mem_2_qos(axi4asink_auto_in_ar_mem_2_qos),
    .auto_in_ar_mem_3_id(axi4asink_auto_in_ar_mem_3_id),
    .auto_in_ar_mem_3_addr(axi4asink_auto_in_ar_mem_3_addr),
    .auto_in_ar_mem_3_len(axi4asink_auto_in_ar_mem_3_len),
    .auto_in_ar_mem_3_size(axi4asink_auto_in_ar_mem_3_size),
    .auto_in_ar_mem_3_burst(axi4asink_auto_in_ar_mem_3_burst),
    .auto_in_ar_mem_3_lock(axi4asink_auto_in_ar_mem_3_lock),
    .auto_in_ar_mem_3_cache(axi4asink_auto_in_ar_mem_3_cache),
    .auto_in_ar_mem_3_prot(axi4asink_auto_in_ar_mem_3_prot),
    .auto_in_ar_mem_3_qos(axi4asink_auto_in_ar_mem_3_qos),
    .auto_in_ar_mem_4_id(axi4asink_auto_in_ar_mem_4_id),
    .auto_in_ar_mem_4_addr(axi4asink_auto_in_ar_mem_4_addr),
    .auto_in_ar_mem_4_len(axi4asink_auto_in_ar_mem_4_len),
    .auto_in_ar_mem_4_size(axi4asink_auto_in_ar_mem_4_size),
    .auto_in_ar_mem_4_burst(axi4asink_auto_in_ar_mem_4_burst),
    .auto_in_ar_mem_4_lock(axi4asink_auto_in_ar_mem_4_lock),
    .auto_in_ar_mem_4_cache(axi4asink_auto_in_ar_mem_4_cache),
    .auto_in_ar_mem_4_prot(axi4asink_auto_in_ar_mem_4_prot),
    .auto_in_ar_mem_4_qos(axi4asink_auto_in_ar_mem_4_qos),
    .auto_in_ar_mem_5_id(axi4asink_auto_in_ar_mem_5_id),
    .auto_in_ar_mem_5_addr(axi4asink_auto_in_ar_mem_5_addr),
    .auto_in_ar_mem_5_len(axi4asink_auto_in_ar_mem_5_len),
    .auto_in_ar_mem_5_size(axi4asink_auto_in_ar_mem_5_size),
    .auto_in_ar_mem_5_burst(axi4asink_auto_in_ar_mem_5_burst),
    .auto_in_ar_mem_5_lock(axi4asink_auto_in_ar_mem_5_lock),
    .auto_in_ar_mem_5_cache(axi4asink_auto_in_ar_mem_5_cache),
    .auto_in_ar_mem_5_prot(axi4asink_auto_in_ar_mem_5_prot),
    .auto_in_ar_mem_5_qos(axi4asink_auto_in_ar_mem_5_qos),
    .auto_in_ar_mem_6_id(axi4asink_auto_in_ar_mem_6_id),
    .auto_in_ar_mem_6_addr(axi4asink_auto_in_ar_mem_6_addr),
    .auto_in_ar_mem_6_len(axi4asink_auto_in_ar_mem_6_len),
    .auto_in_ar_mem_6_size(axi4asink_auto_in_ar_mem_6_size),
    .auto_in_ar_mem_6_burst(axi4asink_auto_in_ar_mem_6_burst),
    .auto_in_ar_mem_6_lock(axi4asink_auto_in_ar_mem_6_lock),
    .auto_in_ar_mem_6_cache(axi4asink_auto_in_ar_mem_6_cache),
    .auto_in_ar_mem_6_prot(axi4asink_auto_in_ar_mem_6_prot),
    .auto_in_ar_mem_6_qos(axi4asink_auto_in_ar_mem_6_qos),
    .auto_in_ar_mem_7_id(axi4asink_auto_in_ar_mem_7_id),
    .auto_in_ar_mem_7_addr(axi4asink_auto_in_ar_mem_7_addr),
    .auto_in_ar_mem_7_len(axi4asink_auto_in_ar_mem_7_len),
    .auto_in_ar_mem_7_size(axi4asink_auto_in_ar_mem_7_size),
    .auto_in_ar_mem_7_burst(axi4asink_auto_in_ar_mem_7_burst),
    .auto_in_ar_mem_7_lock(axi4asink_auto_in_ar_mem_7_lock),
    .auto_in_ar_mem_7_cache(axi4asink_auto_in_ar_mem_7_cache),
    .auto_in_ar_mem_7_prot(axi4asink_auto_in_ar_mem_7_prot),
    .auto_in_ar_mem_7_qos(axi4asink_auto_in_ar_mem_7_qos),
    .auto_in_ar_ridx(axi4asink_auto_in_ar_ridx),
    .auto_in_ar_widx(axi4asink_auto_in_ar_widx),
    .auto_in_ar_safe_ridx_valid(axi4asink_auto_in_ar_safe_ridx_valid),
    .auto_in_ar_safe_widx_valid(axi4asink_auto_in_ar_safe_widx_valid),
    .auto_in_ar_safe_source_reset_n(axi4asink_auto_in_ar_safe_source_reset_n),
    .auto_in_ar_safe_sink_reset_n(axi4asink_auto_in_ar_safe_sink_reset_n),
    .auto_in_r_mem_0_id(axi4asink_auto_in_r_mem_0_id),
    .auto_in_r_mem_0_data(axi4asink_auto_in_r_mem_0_data),
    .auto_in_r_mem_0_resp(axi4asink_auto_in_r_mem_0_resp),
    .auto_in_r_mem_0_last(axi4asink_auto_in_r_mem_0_last),
    .auto_in_r_mem_1_id(axi4asink_auto_in_r_mem_1_id),
    .auto_in_r_mem_1_data(axi4asink_auto_in_r_mem_1_data),
    .auto_in_r_mem_1_resp(axi4asink_auto_in_r_mem_1_resp),
    .auto_in_r_mem_1_last(axi4asink_auto_in_r_mem_1_last),
    .auto_in_r_mem_2_id(axi4asink_auto_in_r_mem_2_id),
    .auto_in_r_mem_2_data(axi4asink_auto_in_r_mem_2_data),
    .auto_in_r_mem_2_resp(axi4asink_auto_in_r_mem_2_resp),
    .auto_in_r_mem_2_last(axi4asink_auto_in_r_mem_2_last),
    .auto_in_r_mem_3_id(axi4asink_auto_in_r_mem_3_id),
    .auto_in_r_mem_3_data(axi4asink_auto_in_r_mem_3_data),
    .auto_in_r_mem_3_resp(axi4asink_auto_in_r_mem_3_resp),
    .auto_in_r_mem_3_last(axi4asink_auto_in_r_mem_3_last),
    .auto_in_r_mem_4_id(axi4asink_auto_in_r_mem_4_id),
    .auto_in_r_mem_4_data(axi4asink_auto_in_r_mem_4_data),
    .auto_in_r_mem_4_resp(axi4asink_auto_in_r_mem_4_resp),
    .auto_in_r_mem_4_last(axi4asink_auto_in_r_mem_4_last),
    .auto_in_r_mem_5_id(axi4asink_auto_in_r_mem_5_id),
    .auto_in_r_mem_5_data(axi4asink_auto_in_r_mem_5_data),
    .auto_in_r_mem_5_resp(axi4asink_auto_in_r_mem_5_resp),
    .auto_in_r_mem_5_last(axi4asink_auto_in_r_mem_5_last),
    .auto_in_r_mem_6_id(axi4asink_auto_in_r_mem_6_id),
    .auto_in_r_mem_6_data(axi4asink_auto_in_r_mem_6_data),
    .auto_in_r_mem_6_resp(axi4asink_auto_in_r_mem_6_resp),
    .auto_in_r_mem_6_last(axi4asink_auto_in_r_mem_6_last),
    .auto_in_r_mem_7_id(axi4asink_auto_in_r_mem_7_id),
    .auto_in_r_mem_7_data(axi4asink_auto_in_r_mem_7_data),
    .auto_in_r_mem_7_resp(axi4asink_auto_in_r_mem_7_resp),
    .auto_in_r_mem_7_last(axi4asink_auto_in_r_mem_7_last),
    .auto_in_r_ridx(axi4asink_auto_in_r_ridx),
    .auto_in_r_widx(axi4asink_auto_in_r_widx),
    .auto_in_r_safe_ridx_valid(axi4asink_auto_in_r_safe_ridx_valid),
    .auto_in_r_safe_widx_valid(axi4asink_auto_in_r_safe_widx_valid),
    .auto_in_r_safe_source_reset_n(axi4asink_auto_in_r_safe_source_reset_n),
    .auto_in_r_safe_sink_reset_n(axi4asink_auto_in_r_safe_sink_reset_n),
    .auto_out_aw_ready(axi4asink_auto_out_aw_ready),
    .auto_out_aw_valid(axi4asink_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4asink_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4asink_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4asink_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4asink_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4asink_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4asink_auto_out_aw_bits_lock),
    .auto_out_aw_bits_prot(axi4asink_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4asink_auto_out_aw_bits_qos),
    .auto_out_w_ready(axi4asink_auto_out_w_ready),
    .auto_out_w_valid(axi4asink_auto_out_w_valid),
    .auto_out_w_bits_data(axi4asink_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4asink_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4asink_auto_out_w_bits_last),
    .auto_out_b_ready(axi4asink_auto_out_b_ready),
    .auto_out_b_valid(axi4asink_auto_out_b_valid),
    .auto_out_b_bits_id(axi4asink_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4asink_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4asink_auto_out_ar_ready),
    .auto_out_ar_valid(axi4asink_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4asink_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4asink_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4asink_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4asink_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4asink_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4asink_auto_out_ar_bits_lock),
    .auto_out_ar_bits_prot(axi4asink_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4asink_auto_out_ar_bits_qos),
    .auto_out_r_ready(axi4asink_auto_out_r_ready),
    .auto_out_r_valid(axi4asink_auto_out_r_valid),
    .auto_out_r_bits_id(axi4asink_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4asink_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4asink_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4asink_auto_out_r_bits_last)
  );
  vc707mig1gb blackbox ( // @[XilinxVC707MIG.scala 53:26:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305220.4]
    .device_temp(blackbox_device_temp),
    .s_axi_rvalid(blackbox_s_axi_rvalid),
    .s_axi_rlast(blackbox_s_axi_rlast),
    .s_axi_rresp(blackbox_s_axi_rresp),
    .s_axi_rdata(blackbox_s_axi_rdata),
    .s_axi_rid(blackbox_s_axi_rid),
    .s_axi_rready(blackbox_s_axi_rready),
    .s_axi_arready(blackbox_s_axi_arready),
    .s_axi_arvalid(blackbox_s_axi_arvalid),
    .s_axi_arqos(blackbox_s_axi_arqos),
    .s_axi_arprot(blackbox_s_axi_arprot),
    .s_axi_arcache(blackbox_s_axi_arcache),
    .s_axi_arlock(blackbox_s_axi_arlock),
    .s_axi_arburst(blackbox_s_axi_arburst),
    .s_axi_arsize(blackbox_s_axi_arsize),
    .s_axi_arlen(blackbox_s_axi_arlen),
    .s_axi_araddr(blackbox_s_axi_araddr),
    .s_axi_arid(blackbox_s_axi_arid),
    .s_axi_bvalid(blackbox_s_axi_bvalid),
    .s_axi_bresp(blackbox_s_axi_bresp),
    .s_axi_bid(blackbox_s_axi_bid),
    .s_axi_bready(blackbox_s_axi_bready),
    .s_axi_wready(blackbox_s_axi_wready),
    .s_axi_wvalid(blackbox_s_axi_wvalid),
    .s_axi_wlast(blackbox_s_axi_wlast),
    .s_axi_wstrb(blackbox_s_axi_wstrb),
    .s_axi_wdata(blackbox_s_axi_wdata),
    .s_axi_awready(blackbox_s_axi_awready),
    .s_axi_awvalid(blackbox_s_axi_awvalid),
    .s_axi_awqos(blackbox_s_axi_awqos),
    .s_axi_awprot(blackbox_s_axi_awprot),
    .s_axi_awcache(blackbox_s_axi_awcache),
    .s_axi_awlock(blackbox_s_axi_awlock),
    .s_axi_awburst(blackbox_s_axi_awburst),
    .s_axi_awsize(blackbox_s_axi_awsize),
    .s_axi_awlen(blackbox_s_axi_awlen),
    .s_axi_awaddr(blackbox_s_axi_awaddr),
    .s_axi_awid(blackbox_s_axi_awid),
    .app_zq_ack(blackbox_app_zq_ack),
    .app_ref_ack(blackbox_app_ref_ack),
    .app_sr_active(blackbox_app_sr_active),
    .app_zq_req(blackbox_app_zq_req),
    .app_ref_req(blackbox_app_ref_req),
    .app_sr_req(blackbox_app_sr_req),
    .sys_rst(blackbox_sys_rst),
    .init_calib_complete(blackbox_init_calib_complete),
    .aresetn(blackbox_aresetn),
    .mmcm_locked(blackbox_mmcm_locked),
    .ui_clk_sync_rst(blackbox_ui_clk_sync_rst),
    .ui_clk(blackbox_ui_clk),
    .sys_clk_i(blackbox_sys_clk_i),
    .ddr3_dqs_p(io_port_ddr3_dqs_p),
    .ddr3_dqs_n(io_port_ddr3_dqs_n),
    .ddr3_dq(io_port_ddr3_dq),
    .ddr3_odt(blackbox_ddr3_odt),
    .ddr3_dm(blackbox_ddr3_dm),
    .ddr3_cs_n(blackbox_ddr3_cs_n),
    .ddr3_cke(blackbox_ddr3_cke),
    .ddr3_ck_n(blackbox_ddr3_ck_n),
    .ddr3_ck_p(blackbox_ddr3_ck_p),
    .ddr3_reset_n(blackbox_ddr3_reset_n),
    .ddr3_we_n(blackbox_ddr3_we_n),
    .ddr3_cas_n(blackbox_ddr3_cas_n),
    .ddr3_ras_n(blackbox_ddr3_ras_n),
    .ddr3_ba(blackbox_ddr3_ba),
    .ddr3_addr(blackbox_ddr3_addr)
  );
  assign axi_async_aw_bits_addr = axi4asink_auto_out_aw_bits_addr; // @[Nodes.scala 333:76:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305208.4 LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign _T_1172 = axi_async_aw_bits_addr - 32'h80000000; // @[XilinxVC707MIG.scala 92:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305310.4]
  assign _T_1173 = $unsigned(_T_1172); // @[XilinxVC707MIG.scala 92:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305311.4]
  assign awaddr = _T_1173[31:0]; // @[XilinxVC707MIG.scala 92:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305312.4]
  assign axi_async_ar_bits_addr = axi4asink_auto_out_ar_bits_addr; // @[Nodes.scala 333:76:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305208.4 LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign _T_1174 = axi_async_ar_bits_addr - 32'h80000000; // @[XilinxVC707MIG.scala 93:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305313.4]
  assign _T_1175 = $unsigned(_T_1174); // @[XilinxVC707MIG.scala 93:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305314.4]
  assign araddr = _T_1175[31:0]; // @[XilinxVC707MIG.scala 93:41:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305315.4]
  assign auto_axi4in_xing_in_aw_ridx = axi4asink_auto_in_aw_ridx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_aw_safe_ridx_valid = axi4asink_auto_in_aw_safe_ridx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_aw_safe_sink_reset_n = axi4asink_auto_in_aw_safe_sink_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_w_ridx = axi4asink_auto_in_w_ridx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_w_safe_ridx_valid = axi4asink_auto_in_w_safe_ridx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_w_safe_sink_reset_n = axi4asink_auto_in_w_safe_sink_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_0_id = axi4asink_auto_in_b_mem_0_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_0_resp = axi4asink_auto_in_b_mem_0_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_1_id = axi4asink_auto_in_b_mem_1_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_1_resp = axi4asink_auto_in_b_mem_1_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_2_id = axi4asink_auto_in_b_mem_2_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_2_resp = axi4asink_auto_in_b_mem_2_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_3_id = axi4asink_auto_in_b_mem_3_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_3_resp = axi4asink_auto_in_b_mem_3_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_4_id = axi4asink_auto_in_b_mem_4_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_4_resp = axi4asink_auto_in_b_mem_4_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_5_id = axi4asink_auto_in_b_mem_5_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_5_resp = axi4asink_auto_in_b_mem_5_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_6_id = axi4asink_auto_in_b_mem_6_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_6_resp = axi4asink_auto_in_b_mem_6_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_7_id = axi4asink_auto_in_b_mem_7_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_mem_7_resp = axi4asink_auto_in_b_mem_7_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_widx = axi4asink_auto_in_b_widx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_safe_widx_valid = axi4asink_auto_in_b_safe_widx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_b_safe_source_reset_n = axi4asink_auto_in_b_safe_source_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_ar_ridx = axi4asink_auto_in_ar_ridx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_ar_safe_ridx_valid = axi4asink_auto_in_ar_safe_ridx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_ar_safe_sink_reset_n = axi4asink_auto_in_ar_safe_sink_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_0_id = axi4asink_auto_in_r_mem_0_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_0_data = axi4asink_auto_in_r_mem_0_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_0_resp = axi4asink_auto_in_r_mem_0_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_0_last = axi4asink_auto_in_r_mem_0_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_1_id = axi4asink_auto_in_r_mem_1_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_1_data = axi4asink_auto_in_r_mem_1_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_1_resp = axi4asink_auto_in_r_mem_1_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_1_last = axi4asink_auto_in_r_mem_1_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_2_id = axi4asink_auto_in_r_mem_2_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_2_data = axi4asink_auto_in_r_mem_2_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_2_resp = axi4asink_auto_in_r_mem_2_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_2_last = axi4asink_auto_in_r_mem_2_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_3_id = axi4asink_auto_in_r_mem_3_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_3_data = axi4asink_auto_in_r_mem_3_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_3_resp = axi4asink_auto_in_r_mem_3_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_3_last = axi4asink_auto_in_r_mem_3_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_4_id = axi4asink_auto_in_r_mem_4_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_4_data = axi4asink_auto_in_r_mem_4_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_4_resp = axi4asink_auto_in_r_mem_4_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_4_last = axi4asink_auto_in_r_mem_4_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_5_id = axi4asink_auto_in_r_mem_5_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_5_data = axi4asink_auto_in_r_mem_5_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_5_resp = axi4asink_auto_in_r_mem_5_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_5_last = axi4asink_auto_in_r_mem_5_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_6_id = axi4asink_auto_in_r_mem_6_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_6_data = axi4asink_auto_in_r_mem_6_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_6_resp = axi4asink_auto_in_r_mem_6_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_6_last = axi4asink_auto_in_r_mem_6_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_7_id = axi4asink_auto_in_r_mem_7_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_7_data = axi4asink_auto_in_r_mem_7_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_7_resp = axi4asink_auto_in_r_mem_7_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_mem_7_last = axi4asink_auto_in_r_mem_7_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_widx = axi4asink_auto_in_r_widx; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_safe_widx_valid = axi4asink_auto_in_r_safe_widx_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign auto_axi4in_xing_in_r_safe_source_reset_n = axi4asink_auto_in_r_safe_source_reset_n; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305217.4]
  assign io_port_ddr3_addr = blackbox_ddr3_addr; // @[XilinxVC707MIG.scala 64:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305290.4]
  assign io_port_ddr3_ba = blackbox_ddr3_ba; // @[XilinxVC707MIG.scala 65:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305291.4]
  assign io_port_ddr3_ras_n = blackbox_ddr3_ras_n; // @[XilinxVC707MIG.scala 66:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305292.4]
  assign io_port_ddr3_cas_n = blackbox_ddr3_cas_n; // @[XilinxVC707MIG.scala 67:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305293.4]
  assign io_port_ddr3_we_n = blackbox_ddr3_we_n; // @[XilinxVC707MIG.scala 68:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305294.4]
  assign io_port_ddr3_reset_n = blackbox_ddr3_reset_n; // @[XilinxVC707MIG.scala 69:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305295.4]
  assign io_port_ddr3_ck_p = blackbox_ddr3_ck_p; // @[XilinxVC707MIG.scala 70:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305296.4]
  assign io_port_ddr3_ck_n = blackbox_ddr3_ck_n; // @[XilinxVC707MIG.scala 71:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305297.4]
  assign io_port_ddr3_cke = blackbox_ddr3_cke; // @[XilinxVC707MIG.scala 72:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305298.4]
  assign io_port_ddr3_cs_n = blackbox_ddr3_cs_n; // @[XilinxVC707MIG.scala 73:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305299.4]
  assign io_port_ddr3_dm = blackbox_ddr3_dm; // @[XilinxVC707MIG.scala 74:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305300.4]
  assign io_port_ddr3_odt = blackbox_ddr3_odt; // @[XilinxVC707MIG.scala 75:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305301.4]
  assign io_port_ui_clk = blackbox_ui_clk; // @[XilinxVC707MIG.scala 81:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305303.4]
  assign io_port_ui_clk_sync_rst = blackbox_ui_clk_sync_rst; // @[XilinxVC707MIG.scala 82:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305304.4]
  assign io_port_mmcm_locked = blackbox_mmcm_locked; // @[XilinxVC707MIG.scala 83:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305305.4]
  assign axi4asink_clock = io_port_ui_clk; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305206.4]
  assign axi4asink_reset = io_port_ui_clk_sync_rst; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305207.4]
  assign axi4asink_auto_in_aw_mem_0_id = auto_axi4in_xing_in_aw_mem_0_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_0_addr = auto_axi4in_xing_in_aw_mem_0_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_0_len = auto_axi4in_xing_in_aw_mem_0_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_0_size = auto_axi4in_xing_in_aw_mem_0_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_0_burst = auto_axi4in_xing_in_aw_mem_0_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_0_lock = auto_axi4in_xing_in_aw_mem_0_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_0_cache = auto_axi4in_xing_in_aw_mem_0_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_0_prot = auto_axi4in_xing_in_aw_mem_0_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_0_qos = auto_axi4in_xing_in_aw_mem_0_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_id = auto_axi4in_xing_in_aw_mem_1_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_addr = auto_axi4in_xing_in_aw_mem_1_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_len = auto_axi4in_xing_in_aw_mem_1_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_size = auto_axi4in_xing_in_aw_mem_1_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_burst = auto_axi4in_xing_in_aw_mem_1_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_lock = auto_axi4in_xing_in_aw_mem_1_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_cache = auto_axi4in_xing_in_aw_mem_1_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_prot = auto_axi4in_xing_in_aw_mem_1_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_1_qos = auto_axi4in_xing_in_aw_mem_1_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_id = auto_axi4in_xing_in_aw_mem_2_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_addr = auto_axi4in_xing_in_aw_mem_2_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_len = auto_axi4in_xing_in_aw_mem_2_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_size = auto_axi4in_xing_in_aw_mem_2_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_burst = auto_axi4in_xing_in_aw_mem_2_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_lock = auto_axi4in_xing_in_aw_mem_2_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_cache = auto_axi4in_xing_in_aw_mem_2_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_prot = auto_axi4in_xing_in_aw_mem_2_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_2_qos = auto_axi4in_xing_in_aw_mem_2_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_id = auto_axi4in_xing_in_aw_mem_3_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_addr = auto_axi4in_xing_in_aw_mem_3_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_len = auto_axi4in_xing_in_aw_mem_3_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_size = auto_axi4in_xing_in_aw_mem_3_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_burst = auto_axi4in_xing_in_aw_mem_3_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_lock = auto_axi4in_xing_in_aw_mem_3_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_cache = auto_axi4in_xing_in_aw_mem_3_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_prot = auto_axi4in_xing_in_aw_mem_3_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_3_qos = auto_axi4in_xing_in_aw_mem_3_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_id = auto_axi4in_xing_in_aw_mem_4_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_addr = auto_axi4in_xing_in_aw_mem_4_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_len = auto_axi4in_xing_in_aw_mem_4_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_size = auto_axi4in_xing_in_aw_mem_4_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_burst = auto_axi4in_xing_in_aw_mem_4_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_lock = auto_axi4in_xing_in_aw_mem_4_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_cache = auto_axi4in_xing_in_aw_mem_4_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_prot = auto_axi4in_xing_in_aw_mem_4_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_4_qos = auto_axi4in_xing_in_aw_mem_4_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_id = auto_axi4in_xing_in_aw_mem_5_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_addr = auto_axi4in_xing_in_aw_mem_5_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_len = auto_axi4in_xing_in_aw_mem_5_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_size = auto_axi4in_xing_in_aw_mem_5_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_burst = auto_axi4in_xing_in_aw_mem_5_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_lock = auto_axi4in_xing_in_aw_mem_5_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_cache = auto_axi4in_xing_in_aw_mem_5_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_prot = auto_axi4in_xing_in_aw_mem_5_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_5_qos = auto_axi4in_xing_in_aw_mem_5_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_id = auto_axi4in_xing_in_aw_mem_6_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_addr = auto_axi4in_xing_in_aw_mem_6_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_len = auto_axi4in_xing_in_aw_mem_6_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_size = auto_axi4in_xing_in_aw_mem_6_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_burst = auto_axi4in_xing_in_aw_mem_6_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_lock = auto_axi4in_xing_in_aw_mem_6_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_cache = auto_axi4in_xing_in_aw_mem_6_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_prot = auto_axi4in_xing_in_aw_mem_6_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_6_qos = auto_axi4in_xing_in_aw_mem_6_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_id = auto_axi4in_xing_in_aw_mem_7_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_addr = auto_axi4in_xing_in_aw_mem_7_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_len = auto_axi4in_xing_in_aw_mem_7_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_size = auto_axi4in_xing_in_aw_mem_7_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_burst = auto_axi4in_xing_in_aw_mem_7_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_lock = auto_axi4in_xing_in_aw_mem_7_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_cache = auto_axi4in_xing_in_aw_mem_7_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_prot = auto_axi4in_xing_in_aw_mem_7_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_mem_7_qos = auto_axi4in_xing_in_aw_mem_7_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_widx = auto_axi4in_xing_in_aw_widx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_safe_widx_valid = auto_axi4in_xing_in_aw_safe_widx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_aw_safe_source_reset_n = auto_axi4in_xing_in_aw_safe_source_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_0_data = auto_axi4in_xing_in_w_mem_0_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_0_strb = auto_axi4in_xing_in_w_mem_0_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_0_last = auto_axi4in_xing_in_w_mem_0_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_1_data = auto_axi4in_xing_in_w_mem_1_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_1_strb = auto_axi4in_xing_in_w_mem_1_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_1_last = auto_axi4in_xing_in_w_mem_1_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_2_data = auto_axi4in_xing_in_w_mem_2_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_2_strb = auto_axi4in_xing_in_w_mem_2_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_2_last = auto_axi4in_xing_in_w_mem_2_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_3_data = auto_axi4in_xing_in_w_mem_3_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_3_strb = auto_axi4in_xing_in_w_mem_3_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_3_last = auto_axi4in_xing_in_w_mem_3_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_4_data = auto_axi4in_xing_in_w_mem_4_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_4_strb = auto_axi4in_xing_in_w_mem_4_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_4_last = auto_axi4in_xing_in_w_mem_4_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_5_data = auto_axi4in_xing_in_w_mem_5_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_5_strb = auto_axi4in_xing_in_w_mem_5_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_5_last = auto_axi4in_xing_in_w_mem_5_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_6_data = auto_axi4in_xing_in_w_mem_6_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_6_strb = auto_axi4in_xing_in_w_mem_6_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_6_last = auto_axi4in_xing_in_w_mem_6_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_7_data = auto_axi4in_xing_in_w_mem_7_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_7_strb = auto_axi4in_xing_in_w_mem_7_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_mem_7_last = auto_axi4in_xing_in_w_mem_7_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_widx = auto_axi4in_xing_in_w_widx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_safe_widx_valid = auto_axi4in_xing_in_w_safe_widx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_w_safe_source_reset_n = auto_axi4in_xing_in_w_safe_source_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_b_ridx = auto_axi4in_xing_in_b_ridx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_b_safe_ridx_valid = auto_axi4in_xing_in_b_safe_ridx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_b_safe_sink_reset_n = auto_axi4in_xing_in_b_safe_sink_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_id = auto_axi4in_xing_in_ar_mem_0_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_addr = auto_axi4in_xing_in_ar_mem_0_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_len = auto_axi4in_xing_in_ar_mem_0_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_size = auto_axi4in_xing_in_ar_mem_0_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_burst = auto_axi4in_xing_in_ar_mem_0_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_lock = auto_axi4in_xing_in_ar_mem_0_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_cache = auto_axi4in_xing_in_ar_mem_0_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_prot = auto_axi4in_xing_in_ar_mem_0_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_0_qos = auto_axi4in_xing_in_ar_mem_0_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_id = auto_axi4in_xing_in_ar_mem_1_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_addr = auto_axi4in_xing_in_ar_mem_1_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_len = auto_axi4in_xing_in_ar_mem_1_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_size = auto_axi4in_xing_in_ar_mem_1_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_burst = auto_axi4in_xing_in_ar_mem_1_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_lock = auto_axi4in_xing_in_ar_mem_1_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_cache = auto_axi4in_xing_in_ar_mem_1_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_prot = auto_axi4in_xing_in_ar_mem_1_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_1_qos = auto_axi4in_xing_in_ar_mem_1_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_id = auto_axi4in_xing_in_ar_mem_2_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_addr = auto_axi4in_xing_in_ar_mem_2_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_len = auto_axi4in_xing_in_ar_mem_2_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_size = auto_axi4in_xing_in_ar_mem_2_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_burst = auto_axi4in_xing_in_ar_mem_2_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_lock = auto_axi4in_xing_in_ar_mem_2_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_cache = auto_axi4in_xing_in_ar_mem_2_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_prot = auto_axi4in_xing_in_ar_mem_2_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_2_qos = auto_axi4in_xing_in_ar_mem_2_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_id = auto_axi4in_xing_in_ar_mem_3_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_addr = auto_axi4in_xing_in_ar_mem_3_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_len = auto_axi4in_xing_in_ar_mem_3_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_size = auto_axi4in_xing_in_ar_mem_3_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_burst = auto_axi4in_xing_in_ar_mem_3_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_lock = auto_axi4in_xing_in_ar_mem_3_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_cache = auto_axi4in_xing_in_ar_mem_3_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_prot = auto_axi4in_xing_in_ar_mem_3_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_3_qos = auto_axi4in_xing_in_ar_mem_3_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_id = auto_axi4in_xing_in_ar_mem_4_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_addr = auto_axi4in_xing_in_ar_mem_4_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_len = auto_axi4in_xing_in_ar_mem_4_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_size = auto_axi4in_xing_in_ar_mem_4_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_burst = auto_axi4in_xing_in_ar_mem_4_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_lock = auto_axi4in_xing_in_ar_mem_4_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_cache = auto_axi4in_xing_in_ar_mem_4_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_prot = auto_axi4in_xing_in_ar_mem_4_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_4_qos = auto_axi4in_xing_in_ar_mem_4_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_id = auto_axi4in_xing_in_ar_mem_5_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_addr = auto_axi4in_xing_in_ar_mem_5_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_len = auto_axi4in_xing_in_ar_mem_5_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_size = auto_axi4in_xing_in_ar_mem_5_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_burst = auto_axi4in_xing_in_ar_mem_5_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_lock = auto_axi4in_xing_in_ar_mem_5_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_cache = auto_axi4in_xing_in_ar_mem_5_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_prot = auto_axi4in_xing_in_ar_mem_5_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_5_qos = auto_axi4in_xing_in_ar_mem_5_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_id = auto_axi4in_xing_in_ar_mem_6_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_addr = auto_axi4in_xing_in_ar_mem_6_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_len = auto_axi4in_xing_in_ar_mem_6_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_size = auto_axi4in_xing_in_ar_mem_6_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_burst = auto_axi4in_xing_in_ar_mem_6_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_lock = auto_axi4in_xing_in_ar_mem_6_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_cache = auto_axi4in_xing_in_ar_mem_6_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_prot = auto_axi4in_xing_in_ar_mem_6_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_6_qos = auto_axi4in_xing_in_ar_mem_6_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_id = auto_axi4in_xing_in_ar_mem_7_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_addr = auto_axi4in_xing_in_ar_mem_7_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_len = auto_axi4in_xing_in_ar_mem_7_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_size = auto_axi4in_xing_in_ar_mem_7_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_burst = auto_axi4in_xing_in_ar_mem_7_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_lock = auto_axi4in_xing_in_ar_mem_7_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_cache = auto_axi4in_xing_in_ar_mem_7_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_prot = auto_axi4in_xing_in_ar_mem_7_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_mem_7_qos = auto_axi4in_xing_in_ar_mem_7_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_widx = auto_axi4in_xing_in_ar_widx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_safe_widx_valid = auto_axi4in_xing_in_ar_safe_widx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_ar_safe_source_reset_n = auto_axi4in_xing_in_ar_safe_source_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_r_ridx = auto_axi4in_xing_in_r_ridx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_r_safe_ridx_valid = auto_axi4in_xing_in_r_safe_ridx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_in_r_safe_sink_reset_n = auto_axi4in_xing_in_r_safe_sink_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305216.4]
  assign axi4asink_auto_out_aw_ready = blackbox_s_axi_awready; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_w_ready = blackbox_s_axi_wready; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_b_valid = blackbox_s_axi_bvalid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_b_bits_id = blackbox_s_axi_bid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_b_bits_resp = blackbox_s_axi_bresp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_ar_ready = blackbox_s_axi_arready; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_r_valid = blackbox_s_axi_rvalid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_r_bits_id = blackbox_s_axi_rid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_r_bits_data = blackbox_s_axi_rdata; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_r_bits_resp = blackbox_s_axi_rresp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign axi4asink_auto_out_r_bits_last = blackbox_s_axi_rlast; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305215.4]
  assign blackbox_s_axi_rready = axi4asink_auto_out_r_ready; // @[XilinxVC707MIG.scala 135:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305347.4]
  assign blackbox_s_axi_arvalid = axi4asink_auto_out_ar_valid; // @[XilinxVC707MIG.scala 131:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305345.4]
  assign blackbox_s_axi_arqos = axi4asink_auto_out_ar_bits_qos; // @[XilinxVC707MIG.scala 130:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305344.4]
  assign blackbox_s_axi_arprot = axi4asink_auto_out_ar_bits_prot; // @[XilinxVC707MIG.scala 129:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305343.4]
  assign blackbox_s_axi_arcache = 4'h3; // @[XilinxVC707MIG.scala 128:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305342.4]
  assign blackbox_s_axi_arlock = axi4asink_auto_out_ar_bits_lock; // @[XilinxVC707MIG.scala 127:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305341.4]
  assign blackbox_s_axi_arburst = axi4asink_auto_out_ar_bits_burst; // @[XilinxVC707MIG.scala 126:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305340.4]
  assign blackbox_s_axi_arsize = axi4asink_auto_out_ar_bits_size; // @[XilinxVC707MIG.scala 125:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305339.4]
  assign blackbox_s_axi_arlen = axi4asink_auto_out_ar_bits_len; // @[XilinxVC707MIG.scala 124:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305338.4]
  assign blackbox_s_axi_araddr = araddr[29:0]; // @[XilinxVC707MIG.scala 123:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305337.4]
  assign blackbox_s_axi_arid = axi4asink_auto_out_ar_bits_id; // @[XilinxVC707MIG.scala 122:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305336.4]
  assign blackbox_s_axi_bready = axi4asink_auto_out_b_ready; // @[XilinxVC707MIG.scala 116:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305332.4]
  assign blackbox_s_axi_wvalid = axi4asink_auto_out_w_valid; // @[XilinxVC707MIG.scala 112:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305330.4]
  assign blackbox_s_axi_wlast = axi4asink_auto_out_w_bits_last; // @[XilinxVC707MIG.scala 111:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305329.4]
  assign blackbox_s_axi_wstrb = axi4asink_auto_out_w_bits_strb; // @[XilinxVC707MIG.scala 110:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305328.4]
  assign blackbox_s_axi_wdata = axi4asink_auto_out_w_bits_data; // @[XilinxVC707MIG.scala 109:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305327.4]
  assign blackbox_s_axi_awvalid = axi4asink_auto_out_aw_valid; // @[XilinxVC707MIG.scala 105:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305325.4]
  assign blackbox_s_axi_awqos = axi4asink_auto_out_aw_bits_qos; // @[XilinxVC707MIG.scala 104:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305324.4]
  assign blackbox_s_axi_awprot = axi4asink_auto_out_aw_bits_prot; // @[XilinxVC707MIG.scala 103:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305323.4]
  assign blackbox_s_axi_awcache = 4'h3; // @[XilinxVC707MIG.scala 102:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305322.4]
  assign blackbox_s_axi_awlock = axi4asink_auto_out_aw_bits_lock; // @[XilinxVC707MIG.scala 101:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305321.4]
  assign blackbox_s_axi_awburst = axi4asink_auto_out_aw_bits_burst; // @[XilinxVC707MIG.scala 100:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305320.4]
  assign blackbox_s_axi_awsize = axi4asink_auto_out_aw_bits_size; // @[XilinxVC707MIG.scala 99:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305319.4]
  assign blackbox_s_axi_awlen = axi4asink_auto_out_aw_bits_len; // @[XilinxVC707MIG.scala 98:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305318.4]
  assign blackbox_s_axi_awaddr = awaddr[29:0]; // @[XilinxVC707MIG.scala 97:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305317.4]
  assign blackbox_s_axi_awid = axi4asink_auto_out_aw_bits_id; // @[XilinxVC707MIG.scala 96:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305316.4]
  assign blackbox_app_zq_req = 1'h0; // @[XilinxVC707MIG.scala 87:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305309.4]
  assign blackbox_app_ref_req = 1'h0; // @[XilinxVC707MIG.scala 86:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305308.4]
  assign blackbox_app_sr_req = 1'h0; // @[XilinxVC707MIG.scala 85:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305307.4]
  assign blackbox_sys_rst = io_port_sys_rst; // @[XilinxVC707MIG.scala 144:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305354.4]
  assign blackbox_aresetn = io_port_aresetn; // @[XilinxVC707MIG.scala 84:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305306.4]
  assign blackbox_sys_clk_i = io_port_sys_clk_i; // @[XilinxVC707MIG.scala 79:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@305302.4]
endmodule
module AsyncQueueSource_5( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306271.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306272.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306273.4]
  output        io_enq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input         io_enq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [3:0]  io_enq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [31:0] io_enq_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [7:0]  io_enq_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [2:0]  io_enq_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [1:0]  io_enq_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input         io_enq_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [3:0]  io_enq_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [2:0]  io_enq_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [3:0]  io_enq_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [31:0] io_async_mem_0_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [7:0]  io_async_mem_0_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_0_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [1:0]  io_async_mem_0_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_mem_0_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_0_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_0_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_0_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [31:0] io_async_mem_1_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [7:0]  io_async_mem_1_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_1_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [1:0]  io_async_mem_1_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_mem_1_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_1_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_1_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_1_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [31:0] io_async_mem_2_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [7:0]  io_async_mem_2_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_2_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [1:0]  io_async_mem_2_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_mem_2_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_2_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_2_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_2_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [31:0] io_async_mem_3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [7:0]  io_async_mem_3_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_3_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [1:0]  io_async_mem_3_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_mem_3_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_3_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_3_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_3_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [31:0] io_async_mem_4_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [7:0]  io_async_mem_4_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_4_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [1:0]  io_async_mem_4_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_mem_4_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_4_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_4_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_4_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [31:0] io_async_mem_5_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [7:0]  io_async_mem_5_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_5_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [1:0]  io_async_mem_5_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_mem_5_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_5_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_5_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_5_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [31:0] io_async_mem_6_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [7:0]  io_async_mem_6_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_6_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [1:0]  io_async_mem_6_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_mem_6_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_6_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_6_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_6_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [31:0] io_async_mem_7_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [7:0]  io_async_mem_7_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_7_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [1:0]  io_async_mem_7_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_mem_7_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_7_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [2:0]  io_async_mem_7_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_mem_7_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input  [3:0]  io_async_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output [3:0]  io_async_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input         io_async_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  output        io_async_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
  input         io_async_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306274.4]
);
  wire  widx_bin_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306282.4]
  wire  widx_bin_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306282.4]
  wire [3:0] widx_bin_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306282.4]
  wire [3:0] widx_bin_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306282.4]
  wire  widx_bin_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306282.4]
  wire  ridx_gray_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306294.4]
  wire  ridx_gray_reset; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306294.4]
  wire [3:0] ridx_gray_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306294.4]
  wire [3:0] ridx_gray_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306294.4]
  wire  ready_reg_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306321.4]
  wire  ready_reg_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306321.4]
  wire  ready_reg_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306321.4]
  wire  ready_reg_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306321.4]
  wire  ready_reg_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306321.4]
  wire  widx_gray_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306330.4]
  wire  widx_gray_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306330.4]
  wire [3:0] widx_gray_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306330.4]
  wire [3:0] widx_gray_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306330.4]
  wire  widx_gray_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306330.4]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306409.4]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306409.4]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306409.4]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306409.4]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306412.4]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306412.4]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306412.4]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306412.4]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306415.4]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306415.4]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306415.4]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306415.4]
  reg [3:0] mem_0_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_0;
  reg [31:0] mem_0_addr; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_1;
  reg [7:0] mem_0_len; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_2;
  reg [2:0] mem_0_size; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_3;
  reg [1:0] mem_0_burst; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_4;
  reg  mem_0_lock; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_5;
  reg [3:0] mem_0_cache; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_6;
  reg [2:0] mem_0_prot; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_7;
  reg [3:0] mem_0_qos; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_8;
  reg [3:0] mem_1_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_9;
  reg [31:0] mem_1_addr; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_10;
  reg [7:0] mem_1_len; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_11;
  reg [2:0] mem_1_size; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_12;
  reg [1:0] mem_1_burst; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_13;
  reg  mem_1_lock; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_14;
  reg [3:0] mem_1_cache; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_15;
  reg [2:0] mem_1_prot; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_16;
  reg [3:0] mem_1_qos; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_17;
  reg [3:0] mem_2_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_18;
  reg [31:0] mem_2_addr; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_19;
  reg [7:0] mem_2_len; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_20;
  reg [2:0] mem_2_size; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_21;
  reg [1:0] mem_2_burst; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_22;
  reg  mem_2_lock; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_23;
  reg [3:0] mem_2_cache; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_24;
  reg [2:0] mem_2_prot; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_25;
  reg [3:0] mem_2_qos; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_26;
  reg [3:0] mem_3_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_27;
  reg [31:0] mem_3_addr; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_28;
  reg [7:0] mem_3_len; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_29;
  reg [2:0] mem_3_size; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_30;
  reg [1:0] mem_3_burst; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_31;
  reg  mem_3_lock; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_32;
  reg [3:0] mem_3_cache; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_33;
  reg [2:0] mem_3_prot; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_34;
  reg [3:0] mem_3_qos; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_35;
  reg [3:0] mem_4_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_36;
  reg [31:0] mem_4_addr; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_37;
  reg [7:0] mem_4_len; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_38;
  reg [2:0] mem_4_size; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_39;
  reg [1:0] mem_4_burst; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_40;
  reg  mem_4_lock; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_41;
  reg [3:0] mem_4_cache; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_42;
  reg [2:0] mem_4_prot; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_43;
  reg [3:0] mem_4_qos; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_44;
  reg [3:0] mem_5_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_45;
  reg [31:0] mem_5_addr; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_46;
  reg [7:0] mem_5_len; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_47;
  reg [2:0] mem_5_size; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_48;
  reg [1:0] mem_5_burst; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_49;
  reg  mem_5_lock; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_50;
  reg [3:0] mem_5_cache; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_51;
  reg [2:0] mem_5_prot; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_52;
  reg [3:0] mem_5_qos; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_53;
  reg [3:0] mem_6_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_54;
  reg [31:0] mem_6_addr; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_55;
  reg [7:0] mem_6_len; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_56;
  reg [2:0] mem_6_size; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_57;
  reg [1:0] mem_6_burst; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_58;
  reg  mem_6_lock; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_59;
  reg [3:0] mem_6_cache; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_60;
  reg [2:0] mem_6_prot; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_61;
  reg [3:0] mem_6_qos; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_62;
  reg [3:0] mem_7_id; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_63;
  reg [31:0] mem_7_addr; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_64;
  reg [7:0] mem_7_len; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_65;
  reg [2:0] mem_7_size; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_66;
  reg [1:0] mem_7_burst; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_67;
  reg  mem_7_lock; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_68;
  reg [3:0] mem_7_cache; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_69;
  reg [2:0] mem_7_prot; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_70;
  reg [3:0] mem_7_qos; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306278.4]
  reg [31:0] _RAND_71;
  wire  _T_64; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306279.4]
  wire  sink_ready; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306276.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306277.4 AsyncQueue.scala 106:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306430.4]
  wire  _T_65; // @[AsyncQueue.scala 77:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306280.4]
  wire [3:0] _GEN_144; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306288.4]
  wire [3:0] _T_69; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306289.4]
  wire [3:0] _T_70; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306290.4]
  wire [2:0] _T_71; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306292.4]
  wire [3:0] _GEN_145; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306293.4]
  wire [3:0] widx; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306293.4]
  wire [3:0] ridx; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306299.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306301.4]
  wire [3:0] _T_73; // @[AsyncQueue.scala 79:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306302.4]
  wire  _T_74; // @[AsyncQueue.scala 79:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306303.4]
  wire [2:0] _T_75; // @[AsyncQueue.scala 81:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306305.4]
  wire  _T_76; // @[AsyncQueue.scala 81:80:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306306.4]
  wire [2:0] _GEN_146; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306307.4]
  wire [2:0] _T_77; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306307.4]
  wire [2:0] index; // @[AsyncQueue.scala 81:64:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306308.4]
  wire  ready_reg_1; // @[AsyncQueue.scala 84:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306327.4]
  wire  _T_82; // @[AsyncQueue.scala 99:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306419.4]
  AsyncResetRegVec_w4_i0 widx_bin ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306282.4]
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_gray ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306294.4]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  AsyncResetRegVec_w1_i0 ready_reg ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306321.4]
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_w4_i0 widx_gray ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306330.4]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306409.4]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306412.4]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306415.4]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign _T_64 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306279.4]
  assign sink_ready = AsyncValidSync_2_io_out; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306276.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306277.4 AsyncQueue.scala 106:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306430.4]
  assign _T_65 = sink_ready == 1'h0; // @[AsyncQueue.scala 77:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306280.4]
  assign _GEN_144 = {{3'd0}, _T_64}; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306288.4]
  assign _T_69 = widx_bin_io_q + _GEN_144; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306289.4]
  assign _T_70 = _T_65 ? 4'h0 : _T_69; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306290.4]
  assign _T_71 = _T_70[3:1]; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306292.4]
  assign _GEN_145 = {{1'd0}, _T_71}; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306293.4]
  assign widx = _T_70 ^ _GEN_145; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306293.4]
  assign ridx = ridx_gray_io_q; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306299.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306301.4]
  assign _T_73 = ridx ^ 4'hc; // @[AsyncQueue.scala 79:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306302.4]
  assign _T_74 = widx != _T_73; // @[AsyncQueue.scala 79:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306303.4]
  assign _T_75 = io_async_widx[2:0]; // @[AsyncQueue.scala 81:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306305.4]
  assign _T_76 = io_async_widx[3]; // @[AsyncQueue.scala 81:80:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306306.4]
  assign _GEN_146 = {{2'd0}, _T_76}; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306307.4]
  assign _T_77 = _GEN_146 << 2; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306307.4]
  assign index = _T_75 ^ _T_77; // @[AsyncQueue.scala 81:64:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306308.4]
  assign ready_reg_1 = ready_reg_io_q; // @[AsyncQueue.scala 84:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306327.4]
  assign _T_82 = io_async_safe_sink_reset_n == 1'h0; // @[AsyncQueue.scala 99:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306419.4]
  assign io_enq_ready = ready_reg_1 & sink_ready; // @[AsyncQueue.scala 85:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306329.4]
  assign io_async_mem_0_id = mem_0_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306345.4]
  assign io_async_mem_0_addr = mem_0_addr; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306344.4]
  assign io_async_mem_0_len = mem_0_len; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306343.4]
  assign io_async_mem_0_size = mem_0_size; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306342.4]
  assign io_async_mem_0_burst = mem_0_burst; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306341.4]
  assign io_async_mem_0_lock = mem_0_lock; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306340.4]
  assign io_async_mem_0_cache = mem_0_cache; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306339.4]
  assign io_async_mem_0_prot = mem_0_prot; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306338.4]
  assign io_async_mem_0_qos = mem_0_qos; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306337.4]
  assign io_async_mem_1_id = mem_1_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306354.4]
  assign io_async_mem_1_addr = mem_1_addr; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306353.4]
  assign io_async_mem_1_len = mem_1_len; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306352.4]
  assign io_async_mem_1_size = mem_1_size; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306351.4]
  assign io_async_mem_1_burst = mem_1_burst; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306350.4]
  assign io_async_mem_1_lock = mem_1_lock; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306349.4]
  assign io_async_mem_1_cache = mem_1_cache; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306348.4]
  assign io_async_mem_1_prot = mem_1_prot; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306347.4]
  assign io_async_mem_1_qos = mem_1_qos; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306346.4]
  assign io_async_mem_2_id = mem_2_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306363.4]
  assign io_async_mem_2_addr = mem_2_addr; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306362.4]
  assign io_async_mem_2_len = mem_2_len; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306361.4]
  assign io_async_mem_2_size = mem_2_size; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306360.4]
  assign io_async_mem_2_burst = mem_2_burst; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306359.4]
  assign io_async_mem_2_lock = mem_2_lock; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306358.4]
  assign io_async_mem_2_cache = mem_2_cache; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306357.4]
  assign io_async_mem_2_prot = mem_2_prot; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306356.4]
  assign io_async_mem_2_qos = mem_2_qos; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306355.4]
  assign io_async_mem_3_id = mem_3_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306372.4]
  assign io_async_mem_3_addr = mem_3_addr; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306371.4]
  assign io_async_mem_3_len = mem_3_len; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306370.4]
  assign io_async_mem_3_size = mem_3_size; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306369.4]
  assign io_async_mem_3_burst = mem_3_burst; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306368.4]
  assign io_async_mem_3_lock = mem_3_lock; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306367.4]
  assign io_async_mem_3_cache = mem_3_cache; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306366.4]
  assign io_async_mem_3_prot = mem_3_prot; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306365.4]
  assign io_async_mem_3_qos = mem_3_qos; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306364.4]
  assign io_async_mem_4_id = mem_4_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306381.4]
  assign io_async_mem_4_addr = mem_4_addr; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306380.4]
  assign io_async_mem_4_len = mem_4_len; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306379.4]
  assign io_async_mem_4_size = mem_4_size; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306378.4]
  assign io_async_mem_4_burst = mem_4_burst; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306377.4]
  assign io_async_mem_4_lock = mem_4_lock; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306376.4]
  assign io_async_mem_4_cache = mem_4_cache; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306375.4]
  assign io_async_mem_4_prot = mem_4_prot; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306374.4]
  assign io_async_mem_4_qos = mem_4_qos; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306373.4]
  assign io_async_mem_5_id = mem_5_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306390.4]
  assign io_async_mem_5_addr = mem_5_addr; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306389.4]
  assign io_async_mem_5_len = mem_5_len; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306388.4]
  assign io_async_mem_5_size = mem_5_size; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306387.4]
  assign io_async_mem_5_burst = mem_5_burst; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306386.4]
  assign io_async_mem_5_lock = mem_5_lock; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306385.4]
  assign io_async_mem_5_cache = mem_5_cache; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306384.4]
  assign io_async_mem_5_prot = mem_5_prot; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306383.4]
  assign io_async_mem_5_qos = mem_5_qos; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306382.4]
  assign io_async_mem_6_id = mem_6_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306399.4]
  assign io_async_mem_6_addr = mem_6_addr; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306398.4]
  assign io_async_mem_6_len = mem_6_len; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306397.4]
  assign io_async_mem_6_size = mem_6_size; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306396.4]
  assign io_async_mem_6_burst = mem_6_burst; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306395.4]
  assign io_async_mem_6_lock = mem_6_lock; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306394.4]
  assign io_async_mem_6_cache = mem_6_cache; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306393.4]
  assign io_async_mem_6_prot = mem_6_prot; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306392.4]
  assign io_async_mem_6_qos = mem_6_qos; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306391.4]
  assign io_async_mem_7_id = mem_7_id; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306408.4]
  assign io_async_mem_7_addr = mem_7_addr; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306407.4]
  assign io_async_mem_7_len = mem_7_len; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306406.4]
  assign io_async_mem_7_size = mem_7_size; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306405.4]
  assign io_async_mem_7_burst = mem_7_burst; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306404.4]
  assign io_async_mem_7_lock = mem_7_lock; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306403.4]
  assign io_async_mem_7_cache = mem_7_cache; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306402.4]
  assign io_async_mem_7_prot = mem_7_prot; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306401.4]
  assign io_async_mem_7_qos = mem_7_qos; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306400.4]
  assign io_async_widx = widx_gray_io_q; // @[AsyncQueue.scala 88:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306336.4]
  assign io_async_safe_widx_valid = AsyncValidSync_io_out; // @[AsyncQueue.scala 103:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306427.4]
  assign io_async_safe_source_reset_n = reset == 1'h0; // @[AsyncQueue.scala 107:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306433.4]
  assign widx_bin_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306284.4]
  assign widx_bin_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306285.4]
  assign widx_bin_io_d = _T_65 ? 4'h0 : _T_69; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306286.4]
  assign widx_bin_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306287.4]
  assign ridx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306296.4]
  assign ridx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306297.4]
  assign ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306298.4]
  assign ready_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306323.4]
  assign ready_reg_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306324.4]
  assign ready_reg_io_d = sink_ready & _T_74; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306325.4]
  assign ready_reg_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306326.4]
  assign widx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306332.4]
  assign widx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306333.4]
  assign widx_gray_io_d = _T_70 ^ _GEN_145; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306334.4]
  assign widx_gray_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306335.4]
  assign AsyncValidSync_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306410.4]
  assign AsyncValidSync_reset = reset | _T_82; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306411.4 AsyncQueue.scala 99:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306421.4]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 102:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306426.4]
  assign AsyncValidSync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306413.4]
  assign AsyncValidSync_1_reset = reset | _T_82; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306414.4 AsyncQueue.scala 100:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306425.4]
  assign AsyncValidSync_1_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 104:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306428.4]
  assign AsyncValidSync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306416.4]
  assign AsyncValidSync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306417.4]
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 105:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@306429.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_id = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_0_addr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_0_len = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_0_size = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_0_burst = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_0_lock = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_0_cache = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_0_prot = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_0_qos = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mem_1_id = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_1_addr = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_1_len = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mem_1_size = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mem_1_burst = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mem_1_lock = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mem_1_cache = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  mem_1_prot = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mem_1_qos = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  mem_2_id = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  mem_2_addr = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  mem_2_len = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  mem_2_size = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_2_burst = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_2_lock = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mem_2_cache = _RAND_24[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_2_prot = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_2_qos = _RAND_26[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_3_id = _RAND_27[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_3_addr = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_3_len = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_3_size = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_3_burst = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mem_3_lock = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  mem_3_cache = _RAND_33[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  mem_3_prot = _RAND_34[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  mem_3_qos = _RAND_35[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  mem_4_id = _RAND_36[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  mem_4_addr = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  mem_4_len = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  mem_4_size = _RAND_39[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  mem_4_burst = _RAND_40[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  mem_4_lock = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  mem_4_cache = _RAND_42[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  mem_4_prot = _RAND_43[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  mem_4_qos = _RAND_44[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  mem_5_id = _RAND_45[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  mem_5_addr = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  mem_5_len = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  mem_5_size = _RAND_48[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  mem_5_burst = _RAND_49[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  mem_5_lock = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  mem_5_cache = _RAND_51[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  mem_5_prot = _RAND_52[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  mem_5_qos = _RAND_53[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  mem_6_id = _RAND_54[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  mem_6_addr = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  mem_6_len = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  mem_6_size = _RAND_57[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  mem_6_burst = _RAND_58[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  mem_6_lock = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  mem_6_cache = _RAND_60[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  mem_6_prot = _RAND_61[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  mem_6_qos = _RAND_62[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  mem_7_id = _RAND_63[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  mem_7_addr = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  mem_7_len = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  mem_7_size = _RAND_66[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  mem_7_burst = _RAND_67[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  mem_7_lock = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  mem_7_cache = _RAND_69[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  mem_7_prot = _RAND_70[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  mem_7_qos = _RAND_71[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_addr <= io_enq_bits_addr;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_len <= io_enq_bits_len;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_size <= io_enq_bits_size;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_burst <= io_enq_bits_burst;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_lock <= io_enq_bits_lock;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_cache <= io_enq_bits_cache;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_prot <= io_enq_bits_prot;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_qos <= io_enq_bits_qos;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_addr <= io_enq_bits_addr;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_len <= io_enq_bits_len;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_size <= io_enq_bits_size;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_burst <= io_enq_bits_burst;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_lock <= io_enq_bits_lock;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_cache <= io_enq_bits_cache;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_prot <= io_enq_bits_prot;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_qos <= io_enq_bits_qos;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_addr <= io_enq_bits_addr;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_len <= io_enq_bits_len;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_size <= io_enq_bits_size;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_burst <= io_enq_bits_burst;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_lock <= io_enq_bits_lock;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_cache <= io_enq_bits_cache;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_prot <= io_enq_bits_prot;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_qos <= io_enq_bits_qos;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_addr <= io_enq_bits_addr;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_len <= io_enq_bits_len;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_size <= io_enq_bits_size;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_burst <= io_enq_bits_burst;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_lock <= io_enq_bits_lock;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_cache <= io_enq_bits_cache;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_prot <= io_enq_bits_prot;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_qos <= io_enq_bits_qos;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_addr <= io_enq_bits_addr;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_len <= io_enq_bits_len;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_size <= io_enq_bits_size;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_burst <= io_enq_bits_burst;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_lock <= io_enq_bits_lock;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_cache <= io_enq_bits_cache;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_prot <= io_enq_bits_prot;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_qos <= io_enq_bits_qos;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_addr <= io_enq_bits_addr;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_len <= io_enq_bits_len;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_size <= io_enq_bits_size;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_burst <= io_enq_bits_burst;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_lock <= io_enq_bits_lock;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_cache <= io_enq_bits_cache;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_prot <= io_enq_bits_prot;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_qos <= io_enq_bits_qos;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_addr <= io_enq_bits_addr;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_len <= io_enq_bits_len;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_size <= io_enq_bits_size;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_burst <= io_enq_bits_burst;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_lock <= io_enq_bits_lock;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_cache <= io_enq_bits_cache;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_prot <= io_enq_bits_prot;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_qos <= io_enq_bits_qos;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_id <= io_enq_bits_id;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_addr <= io_enq_bits_addr;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_len <= io_enq_bits_len;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_size <= io_enq_bits_size;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_burst <= io_enq_bits_burst;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_lock <= io_enq_bits_lock;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_cache <= io_enq_bits_cache;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_prot <= io_enq_bits_prot;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_qos <= io_enq_bits_qos;
      end
    end
  end
endmodule
module AsyncQueueSource_7( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308429.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308430.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308431.4]
  output        io_enq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  input         io_enq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  input  [63:0] io_enq_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  input  [7:0]  io_enq_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  input         io_enq_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [63:0] io_async_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [7:0]  io_async_mem_0_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [63:0] io_async_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [7:0]  io_async_mem_1_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [63:0] io_async_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [7:0]  io_async_mem_2_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [63:0] io_async_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [7:0]  io_async_mem_3_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [63:0] io_async_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [7:0]  io_async_mem_4_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [63:0] io_async_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [7:0]  io_async_mem_5_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [63:0] io_async_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [7:0]  io_async_mem_6_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [63:0] io_async_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [7:0]  io_async_mem_7_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  input  [3:0]  io_async_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output [3:0]  io_async_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  input         io_async_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  output        io_async_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
  input         io_async_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308432.4]
);
  wire  widx_bin_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308440.4]
  wire  widx_bin_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308440.4]
  wire [3:0] widx_bin_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308440.4]
  wire [3:0] widx_bin_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308440.4]
  wire  widx_bin_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308440.4]
  wire  ridx_gray_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308452.4]
  wire  ridx_gray_reset; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308452.4]
  wire [3:0] ridx_gray_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308452.4]
  wire [3:0] ridx_gray_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308452.4]
  wire  ready_reg_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308473.4]
  wire  ready_reg_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308473.4]
  wire  ready_reg_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308473.4]
  wire  ready_reg_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308473.4]
  wire  ready_reg_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308473.4]
  wire  widx_gray_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308482.4]
  wire  widx_gray_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308482.4]
  wire [3:0] widx_gray_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308482.4]
  wire [3:0] widx_gray_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308482.4]
  wire  widx_gray_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308482.4]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308513.4]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308513.4]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308513.4]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308513.4]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308516.4]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308516.4]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308516.4]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308516.4]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308519.4]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308519.4]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308519.4]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308519.4]
  reg [63:0] mem_0_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [63:0] _RAND_0;
  reg [7:0] mem_0_strb; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_1;
  reg  mem_0_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_2;
  reg [63:0] mem_1_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [63:0] _RAND_3;
  reg [7:0] mem_1_strb; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_4;
  reg  mem_1_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_5;
  reg [63:0] mem_2_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [63:0] _RAND_6;
  reg [7:0] mem_2_strb; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_7;
  reg  mem_2_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_8;
  reg [63:0] mem_3_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [63:0] _RAND_9;
  reg [7:0] mem_3_strb; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_10;
  reg  mem_3_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_11;
  reg [63:0] mem_4_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [63:0] _RAND_12;
  reg [7:0] mem_4_strb; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_13;
  reg  mem_4_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_14;
  reg [63:0] mem_5_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [63:0] _RAND_15;
  reg [7:0] mem_5_strb; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_16;
  reg  mem_5_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_17;
  reg [63:0] mem_6_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [63:0] _RAND_18;
  reg [7:0] mem_6_strb; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_19;
  reg  mem_6_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_20;
  reg [63:0] mem_7_data; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [63:0] _RAND_21;
  reg [7:0] mem_7_strb; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_22;
  reg  mem_7_last; // @[AsyncQueue.scala 76:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308436.4]
  reg [31:0] _RAND_23;
  wire  _T_64; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308437.4]
  wire  sink_ready; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308434.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308435.4 AsyncQueue.scala 106:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308534.4]
  wire  _T_65; // @[AsyncQueue.scala 77:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308438.4]
  wire [3:0] _GEN_48; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308446.4]
  wire [3:0] _T_69; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308447.4]
  wire [3:0] _T_70; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308448.4]
  wire [2:0] _T_71; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308450.4]
  wire [3:0] _GEN_49; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308451.4]
  wire [3:0] widx; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308451.4]
  wire [3:0] ridx; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308457.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308459.4]
  wire [3:0] _T_73; // @[AsyncQueue.scala 79:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308460.4]
  wire  _T_74; // @[AsyncQueue.scala 79:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308461.4]
  wire [2:0] _T_75; // @[AsyncQueue.scala 81:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308463.4]
  wire  _T_76; // @[AsyncQueue.scala 81:80:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308464.4]
  wire [2:0] _GEN_50; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308465.4]
  wire [2:0] _T_77; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308465.4]
  wire [2:0] index; // @[AsyncQueue.scala 81:64:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308466.4]
  wire  ready_reg_1; // @[AsyncQueue.scala 84:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308479.4]
  wire  _T_82; // @[AsyncQueue.scala 99:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308523.4]
  AsyncResetRegVec_w4_i0 widx_bin ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308440.4]
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_gray ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308452.4]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  AsyncResetRegVec_w1_i0 ready_reg ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308473.4]
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_w4_i0 widx_gray ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308482.4]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 96:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308513.4]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 97:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308516.4]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 98:30:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308519.4]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign _T_64 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308437.4]
  assign sink_ready = AsyncValidSync_2_io_out; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308434.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308435.4 AsyncQueue.scala 106:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308534.4]
  assign _T_65 = sink_ready == 1'h0; // @[AsyncQueue.scala 77:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308438.4]
  assign _GEN_48 = {{3'd0}, _T_64}; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308446.4]
  assign _T_69 = widx_bin_io_q + _GEN_48; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308447.4]
  assign _T_70 = _T_65 ? 4'h0 : _T_69; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308448.4]
  assign _T_71 = _T_70[3:1]; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308450.4]
  assign _GEN_49 = {{1'd0}, _T_71}; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308451.4]
  assign widx = _T_70 ^ _GEN_49; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308451.4]
  assign ridx = ridx_gray_io_q; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308457.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308459.4]
  assign _T_73 = ridx ^ 4'hc; // @[AsyncQueue.scala 79:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308460.4]
  assign _T_74 = widx != _T_73; // @[AsyncQueue.scala 79:34:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308461.4]
  assign _T_75 = io_async_widx[2:0]; // @[AsyncQueue.scala 81:52:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308463.4]
  assign _T_76 = io_async_widx[3]; // @[AsyncQueue.scala 81:80:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308464.4]
  assign _GEN_50 = {{2'd0}, _T_76}; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308465.4]
  assign _T_77 = _GEN_50 << 2; // @[AsyncQueue.scala 81:93:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308465.4]
  assign index = _T_75 ^ _T_77; // @[AsyncQueue.scala 81:64:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308466.4]
  assign ready_reg_1 = ready_reg_io_q; // @[AsyncQueue.scala 84:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308479.4]
  assign _T_82 = io_async_safe_sink_reset_n == 1'h0; // @[AsyncQueue.scala 99:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308523.4]
  assign io_enq_ready = ready_reg_1 & sink_ready; // @[AsyncQueue.scala 85:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308481.4]
  assign io_async_mem_0_data = mem_0_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308491.4]
  assign io_async_mem_0_strb = mem_0_strb; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308490.4]
  assign io_async_mem_0_last = mem_0_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308489.4]
  assign io_async_mem_1_data = mem_1_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308494.4]
  assign io_async_mem_1_strb = mem_1_strb; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308493.4]
  assign io_async_mem_1_last = mem_1_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308492.4]
  assign io_async_mem_2_data = mem_2_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308497.4]
  assign io_async_mem_2_strb = mem_2_strb; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308496.4]
  assign io_async_mem_2_last = mem_2_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308495.4]
  assign io_async_mem_3_data = mem_3_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308500.4]
  assign io_async_mem_3_strb = mem_3_strb; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308499.4]
  assign io_async_mem_3_last = mem_3_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308498.4]
  assign io_async_mem_4_data = mem_4_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308503.4]
  assign io_async_mem_4_strb = mem_4_strb; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308502.4]
  assign io_async_mem_4_last = mem_4_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308501.4]
  assign io_async_mem_5_data = mem_5_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308506.4]
  assign io_async_mem_5_strb = mem_5_strb; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308505.4]
  assign io_async_mem_5_last = mem_5_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308504.4]
  assign io_async_mem_6_data = mem_6_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308509.4]
  assign io_async_mem_6_strb = mem_6_strb; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308508.4]
  assign io_async_mem_6_last = mem_6_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308507.4]
  assign io_async_mem_7_data = mem_7_data; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308512.4]
  assign io_async_mem_7_strb = mem_7_strb; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308511.4]
  assign io_async_mem_7_last = mem_7_last; // @[AsyncQueue.scala 92:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308510.4]
  assign io_async_widx = widx_gray_io_q; // @[AsyncQueue.scala 88:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308488.4]
  assign io_async_safe_widx_valid = AsyncValidSync_io_out; // @[AsyncQueue.scala 103:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308531.4]
  assign io_async_safe_source_reset_n = reset == 1'h0; // @[AsyncQueue.scala 107:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308537.4]
  assign widx_bin_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308442.4]
  assign widx_bin_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308443.4]
  assign widx_bin_io_d = _T_65 ? 4'h0 : _T_69; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308444.4]
  assign widx_bin_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308445.4]
  assign ridx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308454.4]
  assign ridx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308455.4]
  assign ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308456.4]
  assign ready_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308475.4]
  assign ready_reg_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308476.4]
  assign ready_reg_io_d = sink_ready & _T_74; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308477.4]
  assign ready_reg_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308478.4]
  assign widx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308484.4]
  assign widx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308485.4]
  assign widx_gray_io_d = _T_70 ^ _GEN_49; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308486.4]
  assign widx_gray_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308487.4]
  assign AsyncValidSync_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308514.4]
  assign AsyncValidSync_reset = reset | _T_82; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308515.4 AsyncQueue.scala 99:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308525.4]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 102:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308530.4]
  assign AsyncValidSync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308517.4]
  assign AsyncValidSync_1_reset = reset | _T_82; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308518.4 AsyncQueue.scala 100:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308529.4]
  assign AsyncValidSync_1_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 104:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308532.4]
  assign AsyncValidSync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308520.4]
  assign AsyncValidSync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308521.4]
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 105:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308533.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mem_0_data = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_0_strb = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_0_last = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  mem_1_data = _RAND_3[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_1_strb = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_1_last = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{`RANDOM}};
  mem_2_data = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_2_strb = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_2_last = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  mem_3_data = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_3_strb = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_3_last = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  mem_4_data = _RAND_12[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mem_4_strb = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mem_4_last = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  mem_5_data = _RAND_15[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  mem_5_strb = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mem_5_last = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  mem_6_data = _RAND_18[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  mem_6_strb = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  mem_6_last = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  mem_7_data = _RAND_21[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_7_strb = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_7_last = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_strb <= io_enq_bits_strb;
      end
    end
    if (_T_64) begin
      if (3'h0 == index) begin
        mem_0_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_strb <= io_enq_bits_strb;
      end
    end
    if (_T_64) begin
      if (3'h1 == index) begin
        mem_1_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_strb <= io_enq_bits_strb;
      end
    end
    if (_T_64) begin
      if (3'h2 == index) begin
        mem_2_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_strb <= io_enq_bits_strb;
      end
    end
    if (_T_64) begin
      if (3'h3 == index) begin
        mem_3_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_strb <= io_enq_bits_strb;
      end
    end
    if (_T_64) begin
      if (3'h4 == index) begin
        mem_4_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_strb <= io_enq_bits_strb;
      end
    end
    if (_T_64) begin
      if (3'h5 == index) begin
        mem_5_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_strb <= io_enq_bits_strb;
      end
    end
    if (_T_64) begin
      if (3'h6 == index) begin
        mem_6_last <= io_enq_bits_last;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_data <= io_enq_bits_data;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_strb <= io_enq_bits_strb;
      end
    end
    if (_T_64) begin
      if (3'h7 == index) begin
        mem_7_last <= io_enq_bits_last;
      end
    end
  end
endmodule
module SynchronizerShiftReg_w71_d1( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308955.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308956.4]
  input  [70:0] io_d, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308958.4]
  output [70:0] io_q // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308958.4]
);
  reg [70:0] sync_0; // @[ShiftReg.scala 114:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308963.4]
  reg [95:0] _RAND_0;
  assign io_q = sync_0; // @[ShiftReg.scala 123:8:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@308965.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  sync_0 = _RAND_0[70:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    sync_0 <= io_d;
  end
endmodule
module AsyncQueueSink_6( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309497.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309498.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309499.4]
  input         io_deq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  output        io_deq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  output [3:0]  io_deq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  output [63:0] io_deq_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  output [1:0]  io_deq_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  output        io_deq_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [63:0] io_async_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [1:0]  io_async_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [63:0] io_async_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [1:0]  io_async_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [63:0] io_async_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [1:0]  io_async_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [63:0] io_async_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [1:0]  io_async_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [63:0] io_async_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [1:0]  io_async_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [63:0] io_async_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [1:0]  io_async_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [63:0] io_async_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [1:0]  io_async_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [63:0] io_async_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [1:0]  io_async_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  output [3:0]  io_async_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input  [3:0]  io_async_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  output        io_async_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  input         io_async_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
  output        io_async_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309500.4]
);
  wire  ridx_bin_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309507.4]
  wire  ridx_bin_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309507.4]
  wire [3:0] ridx_bin_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309507.4]
  wire [3:0] ridx_bin_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309507.4]
  wire  ridx_bin_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309507.4]
  wire  widx_gray_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309519.4]
  wire  widx_gray_reset; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309519.4]
  wire [3:0] widx_gray_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309519.4]
  wire [3:0] widx_gray_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309519.4]
  wire  deq_bits_reg_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309534.4]
  wire [70:0] deq_bits_reg_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309534.4]
  wire [70:0] deq_bits_reg_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309534.4]
  wire  valid_reg_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309559.4]
  wire  valid_reg_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309559.4]
  wire  valid_reg_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309559.4]
  wire  valid_reg_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309559.4]
  wire  valid_reg_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309559.4]
  wire  ridx_gray_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309568.4]
  wire  ridx_gray_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309568.4]
  wire [3:0] ridx_gray_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309568.4]
  wire [3:0] ridx_gray_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309568.4]
  wire  ridx_gray_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309568.4]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309575.4]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309575.4]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309575.4]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309575.4]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309578.4]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309578.4]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309578.4]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309578.4]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309581.4]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309581.4]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309581.4]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309581.4]
  wire  AsyncResetRegVec_w1_i0_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309610.4]
  wire  AsyncResetRegVec_w1_i0_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309610.4]
  wire  AsyncResetRegVec_w1_i0_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309610.4]
  wire  AsyncResetRegVec_w1_i0_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309610.4]
  wire  AsyncResetRegVec_w1_i0_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309610.4]
  wire  _T_86; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309504.4]
  wire  source_ready; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309502.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309503.4 AsyncQueue.scala 164:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309596.4]
  wire  _T_87; // @[AsyncQueue.scala 130:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309505.4]
  wire [3:0] _GEN_32; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309513.4]
  wire [3:0] _T_91; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309514.4]
  wire [3:0] _T_92; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309515.4]
  wire [2:0] _T_93; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309517.4]
  wire [3:0] _GEN_33; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309518.4]
  wire [3:0] ridx; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309518.4]
  wire [3:0] widx; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309524.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309526.4]
  wire  _T_95; // @[AsyncQueue.scala 132:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309527.4]
  wire  valid; // @[AsyncQueue.scala 132:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309528.4]
  wire [2:0] _T_96; // @[AsyncQueue.scala 138:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309529.4]
  wire  _T_97; // @[AsyncQueue.scala 138:62:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309530.4]
  wire [2:0] _GEN_34; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309531.4]
  wire [2:0] _T_98; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309531.4]
  wire [2:0] index; // @[AsyncQueue.scala 138:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309532.4]
  wire [3:0] _GEN_4; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [63:0] _GEN_5; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [1:0] _GEN_6; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire  _GEN_7; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [3:0] _GEN_8; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [63:0] _GEN_9; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [1:0] _GEN_10; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire  _GEN_11; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [3:0] _GEN_12; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [63:0] _GEN_13; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [1:0] _GEN_14; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire  _GEN_15; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [3:0] _GEN_16; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [63:0] _GEN_17; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [1:0] _GEN_18; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire  _GEN_19; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [3:0] _GEN_20; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [63:0] _GEN_21; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [1:0] _GEN_22; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire  _GEN_23; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [3:0] _GEN_24; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [63:0] _GEN_25; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [1:0] _GEN_26; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire  _GEN_27; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [3:0] _GEN_28; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [63:0] _GEN_29; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [1:0] _GEN_30; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire  _GEN_31; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [3:0] deq_bits_nxt_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [63:0] deq_bits_nxt_data; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [1:0] deq_bits_nxt_resp; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire  deq_bits_nxt_last; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  wire [2:0] _T_100; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309538.4]
  wire [67:0] _T_101; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309539.4]
  wire [70:0] _T_106; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309544.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309546.4]
  wire  valid_reg_1; // @[AsyncQueue.scala 147:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309565.4]
  wire  _T_113; // @[AsyncQueue.scala 157:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309585.4]
  AsyncResetRegVec_w4_i0 ridx_bin ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309507.4]
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_gray ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309519.4]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  SynchronizerShiftReg_w71_d1 deq_bits_reg ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309534.4]
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q)
  );
  AsyncResetRegVec_w1_i0 valid_reg ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309559.4]
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_w4_i0 ridx_gray ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309568.4]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309575.4]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309578.4]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309581.4]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309610.4]
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q),
    .io_en(AsyncResetRegVec_w1_i0_io_en)
  );
  assign _T_86 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309504.4]
  assign source_ready = AsyncValidSync_2_io_out; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309502.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309503.4 AsyncQueue.scala 164:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309596.4]
  assign _T_87 = source_ready == 1'h0; // @[AsyncQueue.scala 130:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309505.4]
  assign _GEN_32 = {{3'd0}, _T_86}; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309513.4]
  assign _T_91 = ridx_bin_io_q + _GEN_32; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309514.4]
  assign _T_92 = _T_87 ? 4'h0 : _T_91; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309515.4]
  assign _T_93 = _T_92[3:1]; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309517.4]
  assign _GEN_33 = {{1'd0}, _T_93}; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309518.4]
  assign ridx = _T_92 ^ _GEN_33; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309518.4]
  assign widx = widx_gray_io_q; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309524.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309526.4]
  assign _T_95 = ridx != widx; // @[AsyncQueue.scala 132:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309527.4]
  assign valid = source_ready & _T_95; // @[AsyncQueue.scala 132:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309528.4]
  assign _T_96 = ridx[2:0]; // @[AsyncQueue.scala 138:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309529.4]
  assign _T_97 = ridx[3]; // @[AsyncQueue.scala 138:62:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309530.4]
  assign _GEN_34 = {{2'd0}, _T_97}; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309531.4]
  assign _T_98 = _GEN_34 << 2; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309531.4]
  assign index = _T_96 ^ _T_98; // @[AsyncQueue.scala 138:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309532.4]
  assign _GEN_4 = 3'h1 == index ? io_async_mem_1_id : io_async_mem_0_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_5 = 3'h1 == index ? io_async_mem_1_data : io_async_mem_0_data; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_6 = 3'h1 == index ? io_async_mem_1_resp : io_async_mem_0_resp; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_7 = 3'h1 == index ? io_async_mem_1_last : io_async_mem_0_last; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_8 = 3'h2 == index ? io_async_mem_2_id : _GEN_4; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_9 = 3'h2 == index ? io_async_mem_2_data : _GEN_5; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_10 = 3'h2 == index ? io_async_mem_2_resp : _GEN_6; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_11 = 3'h2 == index ? io_async_mem_2_last : _GEN_7; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_12 = 3'h3 == index ? io_async_mem_3_id : _GEN_8; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_13 = 3'h3 == index ? io_async_mem_3_data : _GEN_9; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_14 = 3'h3 == index ? io_async_mem_3_resp : _GEN_10; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_15 = 3'h3 == index ? io_async_mem_3_last : _GEN_11; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_16 = 3'h4 == index ? io_async_mem_4_id : _GEN_12; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_17 = 3'h4 == index ? io_async_mem_4_data : _GEN_13; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_18 = 3'h4 == index ? io_async_mem_4_resp : _GEN_14; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_19 = 3'h4 == index ? io_async_mem_4_last : _GEN_15; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_20 = 3'h5 == index ? io_async_mem_5_id : _GEN_16; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_21 = 3'h5 == index ? io_async_mem_5_data : _GEN_17; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_22 = 3'h5 == index ? io_async_mem_5_resp : _GEN_18; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_23 = 3'h5 == index ? io_async_mem_5_last : _GEN_19; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_24 = 3'h6 == index ? io_async_mem_6_id : _GEN_20; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_25 = 3'h6 == index ? io_async_mem_6_data : _GEN_21; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_26 = 3'h6 == index ? io_async_mem_6_resp : _GEN_22; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_27 = 3'h6 == index ? io_async_mem_6_last : _GEN_23; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_28 = 3'h7 == index ? io_async_mem_7_id : _GEN_24; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_29 = 3'h7 == index ? io_async_mem_7_data : _GEN_25; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_30 = 3'h7 == index ? io_async_mem_7_resp : _GEN_26; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _GEN_31 = 3'h7 == index ? io_async_mem_7_last : _GEN_27; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign deq_bits_nxt_id = valid ? _GEN_28 : io_deq_bits_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign deq_bits_nxt_data = valid ? _GEN_29 : io_deq_bits_data; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign deq_bits_nxt_resp = valid ? _GEN_30 : io_deq_bits_resp; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign deq_bits_nxt_last = valid ? _GEN_31 : io_deq_bits_last; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309533.4]
  assign _T_100 = {deq_bits_nxt_resp,deq_bits_nxt_last}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309538.4]
  assign _T_101 = {deq_bits_nxt_id,deq_bits_nxt_data}; // @[ShiftReg.scala 49:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309539.4]
  assign _T_106 = deq_bits_reg_io_q; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309544.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309546.4]
  assign valid_reg_1 = valid_reg_io_q; // @[AsyncQueue.scala 147:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309565.4]
  assign _T_113 = io_async_safe_source_reset_n == 1'h0; // @[AsyncQueue.scala 157:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309585.4]
  assign io_deq_valid = valid_reg_1 & source_ready; // @[AsyncQueue.scala 148:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309567.4]
  assign io_deq_bits_id = _T_106[70:67]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309558.4]
  assign io_deq_bits_data = _T_106[66:3]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309557.4]
  assign io_deq_bits_resp = _T_106[2:1]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309556.4]
  assign io_deq_bits_last = _T_106[0]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309555.4]
  assign io_async_ridx = ridx_gray_io_q; // @[AsyncQueue.scala 151:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309574.4]
  assign io_async_safe_ridx_valid = AsyncValidSync_io_out; // @[AsyncQueue.scala 161:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309593.4]
  assign io_async_safe_sink_reset_n = reset == 1'h0; // @[AsyncQueue.scala 165:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309599.4]
  assign ridx_bin_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309509.4]
  assign ridx_bin_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309510.4]
  assign ridx_bin_io_d = _T_87 ? 4'h0 : _T_91; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309511.4]
  assign ridx_bin_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309512.4]
  assign widx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309521.4]
  assign widx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309522.4]
  assign widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309523.4]
  assign deq_bits_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309536.4]
  assign deq_bits_reg_io_d = {_T_101,_T_100}; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309541.4]
  assign valid_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309561.4]
  assign valid_reg_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309562.4]
  assign valid_reg_io_d = source_ready & _T_95; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309563.4]
  assign valid_reg_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309564.4]
  assign ridx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309570.4]
  assign ridx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309571.4]
  assign ridx_gray_io_d = _T_92 ^ _GEN_33; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309572.4]
  assign ridx_gray_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309573.4]
  assign AsyncValidSync_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309576.4]
  assign AsyncValidSync_reset = reset | _T_113; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309577.4 AsyncQueue.scala 157:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309587.4]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 160:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309592.4]
  assign AsyncValidSync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309579.4]
  assign AsyncValidSync_1_reset = reset | _T_113; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309580.4 AsyncQueue.scala 158:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309591.4]
  assign AsyncValidSync_1_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 162:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309594.4]
  assign AsyncValidSync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309582.4]
  assign AsyncValidSync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309583.4]
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 163:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309595.4]
  assign AsyncResetRegVec_w1_i0_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309612.4]
  assign AsyncResetRegVec_w1_i0_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309613.4]
  assign AsyncResetRegVec_w1_i0_io_d = io_async_widx == io_async_ridx; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309614.4]
  assign AsyncResetRegVec_w1_i0_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@309615.4]
endmodule
module SynchronizerShiftReg_w6_d1( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310033.2]
  input        clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310034.4]
  input  [5:0] io_d, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310036.4]
  output [5:0] io_q // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310036.4]
);
  reg [5:0] sync_0; // @[ShiftReg.scala 114:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310041.4]
  reg [31:0] _RAND_0;
  assign io_q = sync_0; // @[ShiftReg.scala 123:8:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310043.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_0 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    sync_0 <= io_d;
  end
endmodule
module AsyncQueueSink_7( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310575.2]
  input        clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310576.4]
  input        reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310577.4]
  input        io_deq_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  output       io_deq_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  output [3:0] io_deq_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  output [1:0] io_deq_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [1:0] io_async_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [1:0] io_async_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [1:0] io_async_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [1:0] io_async_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [1:0] io_async_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [1:0] io_async_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [1:0] io_async_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [1:0] io_async_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  output [3:0] io_async_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input  [3:0] io_async_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  output       io_async_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input        io_async_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  input        io_async_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
  output       io_async_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310578.4]
);
  wire  ridx_bin_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310585.4]
  wire  ridx_bin_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310585.4]
  wire [3:0] ridx_bin_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310585.4]
  wire [3:0] ridx_bin_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310585.4]
  wire  ridx_bin_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310585.4]
  wire  widx_gray_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310597.4]
  wire  widx_gray_reset; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310597.4]
  wire [3:0] widx_gray_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310597.4]
  wire [3:0] widx_gray_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310597.4]
  wire  deq_bits_reg_clock; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310612.4]
  wire [5:0] deq_bits_reg_io_d; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310612.4]
  wire [5:0] deq_bits_reg_io_q; // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310612.4]
  wire  valid_reg_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310629.4]
  wire  valid_reg_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310629.4]
  wire  valid_reg_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310629.4]
  wire  valid_reg_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310629.4]
  wire  valid_reg_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310629.4]
  wire  ridx_gray_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310638.4]
  wire  ridx_gray_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310638.4]
  wire [3:0] ridx_gray_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310638.4]
  wire [3:0] ridx_gray_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310638.4]
  wire  ridx_gray_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310638.4]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310645.4]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310645.4]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310645.4]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310645.4]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310648.4]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310648.4]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310648.4]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310648.4]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310651.4]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310651.4]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310651.4]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310651.4]
  wire  AsyncResetRegVec_w1_i0_clock; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310680.4]
  wire  AsyncResetRegVec_w1_i0_reset; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310680.4]
  wire  AsyncResetRegVec_w1_i0_io_d; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310680.4]
  wire  AsyncResetRegVec_w1_i0_io_q; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310680.4]
  wire  AsyncResetRegVec_w1_i0_io_en; // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310680.4]
  wire  _T_86; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310582.4]
  wire  source_ready; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310580.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310581.4 AsyncQueue.scala 164:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310666.4]
  wire  _T_87; // @[AsyncQueue.scala 130:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310583.4]
  wire [3:0] _GEN_16; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310591.4]
  wire [3:0] _T_91; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310592.4]
  wire [3:0] _T_92; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310593.4]
  wire [2:0] _T_93; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310595.4]
  wire [3:0] _GEN_17; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310596.4]
  wire [3:0] ridx; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310596.4]
  wire [3:0] widx; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310602.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310604.4]
  wire  _T_95; // @[AsyncQueue.scala 132:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310605.4]
  wire  valid; // @[AsyncQueue.scala 132:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310606.4]
  wire [2:0] _T_96; // @[AsyncQueue.scala 138:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310607.4]
  wire  _T_97; // @[AsyncQueue.scala 138:62:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310608.4]
  wire [2:0] _GEN_18; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310609.4]
  wire [2:0] _T_98; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310609.4]
  wire [2:0] index; // @[AsyncQueue.scala 138:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310610.4]
  wire [3:0] _GEN_2; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [1:0] _GEN_3; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [3:0] _GEN_4; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [1:0] _GEN_5; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [3:0] _GEN_6; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [1:0] _GEN_7; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [3:0] _GEN_8; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [1:0] _GEN_9; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [3:0] _GEN_10; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [1:0] _GEN_11; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [3:0] _GEN_12; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [1:0] _GEN_13; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [3:0] _GEN_14; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [1:0] _GEN_15; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [3:0] deq_bits_nxt_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [1:0] deq_bits_nxt_resp; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  wire [5:0] _T_104; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310620.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310622.4]
  wire  valid_reg_1; // @[AsyncQueue.scala 147:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310635.4]
  wire  _T_109; // @[AsyncQueue.scala 157:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310655.4]
  AsyncResetRegVec_w4_i0 ridx_bin ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310585.4]
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_gray ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310597.4]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  SynchronizerShiftReg_w6_d1 deq_bits_reg ( // @[ShiftReg.scala 47:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310612.4]
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q)
  );
  AsyncResetRegVec_w1_i0 valid_reg ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310629.4]
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_w4_i0 ridx_gray ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310638.4]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 154:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310645.4]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 155:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310648.4]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 156:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310651.4]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 ( // @[AsyncResetReg.scala 97:21:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310680.4]
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q),
    .io_en(AsyncResetRegVec_w1_i0_io_en)
  );
  assign _T_86 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310582.4]
  assign source_ready = AsyncValidSync_2_io_out; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310580.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310581.4 AsyncQueue.scala 164:18:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310666.4]
  assign _T_87 = source_ready == 1'h0; // @[AsyncQueue.scala 130:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310583.4]
  assign _GEN_16 = {{3'd0}, _T_86}; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310591.4]
  assign _T_91 = ridx_bin_io_q + _GEN_16; // @[AsyncQueue.scala 53:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310592.4]
  assign _T_92 = _T_87 ? 4'h0 : _T_91; // @[AsyncQueue.scala 53:23:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310593.4]
  assign _T_93 = _T_92[3:1]; // @[AsyncQueue.scala 54:32:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310595.4]
  assign _GEN_17 = {{1'd0}, _T_93}; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310596.4]
  assign ridx = _T_92 ^ _GEN_17; // @[AsyncQueue.scala 54:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310596.4]
  assign widx = widx_gray_io_q; // @[ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310602.4 ShiftReg.scala 50:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310604.4]
  assign _T_95 = ridx != widx; // @[AsyncQueue.scala 132:36:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310605.4]
  assign valid = source_ready & _T_95; // @[AsyncQueue.scala 132:28:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310606.4]
  assign _T_96 = ridx[2:0]; // @[AsyncQueue.scala 138:43:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310607.4]
  assign _T_97 = ridx[3]; // @[AsyncQueue.scala 138:62:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310608.4]
  assign _GEN_18 = {{2'd0}, _T_97}; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310609.4]
  assign _T_98 = _GEN_18 << 2; // @[AsyncQueue.scala 138:75:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310609.4]
  assign index = _T_96 ^ _T_98; // @[AsyncQueue.scala 138:55:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310610.4]
  assign _GEN_2 = 3'h1 == index ? io_async_mem_1_id : io_async_mem_0_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_3 = 3'h1 == index ? io_async_mem_1_resp : io_async_mem_0_resp; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_4 = 3'h2 == index ? io_async_mem_2_id : _GEN_2; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_5 = 3'h2 == index ? io_async_mem_2_resp : _GEN_3; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_6 = 3'h3 == index ? io_async_mem_3_id : _GEN_4; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_7 = 3'h3 == index ? io_async_mem_3_resp : _GEN_5; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_8 = 3'h4 == index ? io_async_mem_4_id : _GEN_6; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_9 = 3'h4 == index ? io_async_mem_4_resp : _GEN_7; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_10 = 3'h5 == index ? io_async_mem_5_id : _GEN_8; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_11 = 3'h5 == index ? io_async_mem_5_resp : _GEN_9; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_12 = 3'h6 == index ? io_async_mem_6_id : _GEN_10; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_13 = 3'h6 == index ? io_async_mem_6_resp : _GEN_11; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_14 = 3'h7 == index ? io_async_mem_7_id : _GEN_12; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _GEN_15 = 3'h7 == index ? io_async_mem_7_resp : _GEN_13; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign deq_bits_nxt_id = valid ? _GEN_14 : io_deq_bits_id; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign deq_bits_nxt_resp = valid ? _GEN_15 : io_deq_bits_resp; // @[AsyncQueue.scala 144:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310611.4]
  assign _T_104 = deq_bits_reg_io_q; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310620.4 :sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310622.4]
  assign valid_reg_1 = valid_reg_io_q; // @[AsyncQueue.scala 147:59:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310635.4]
  assign _T_109 = io_async_safe_source_reset_n == 1'h0; // @[AsyncQueue.scala 157:44:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310655.4]
  assign io_deq_valid = valid_reg_1 & source_ready; // @[AsyncQueue.scala 148:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310637.4]
  assign io_deq_bits_id = _T_104[5:2]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310628.4]
  assign io_deq_bits_resp = _T_104[1:0]; // @[AsyncQueue.scala 145:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310627.4]
  assign io_async_ridx = ridx_gray_io_q; // @[AsyncQueue.scala 151:17:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310644.4]
  assign io_async_safe_ridx_valid = AsyncValidSync_io_out; // @[AsyncQueue.scala 161:20:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310663.4]
  assign io_async_safe_sink_reset_n = reset == 1'h0; // @[AsyncQueue.scala 165:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310669.4]
  assign ridx_bin_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310587.4]
  assign ridx_bin_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310588.4]
  assign ridx_bin_io_d = _T_87 ? 4'h0 : _T_91; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310589.4]
  assign ridx_bin_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310590.4]
  assign widx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310599.4]
  assign widx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310600.4]
  assign widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310601.4]
  assign deq_bits_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310614.4]
  assign deq_bits_reg_io_d = {deq_bits_nxt_id,deq_bits_nxt_resp}; // @[ShiftReg.scala 49:16:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310617.4]
  assign valid_reg_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310631.4]
  assign valid_reg_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310632.4]
  assign valid_reg_io_d = source_ready & _T_95; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310633.4]
  assign valid_reg_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310634.4]
  assign ridx_gray_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310640.4]
  assign ridx_gray_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310641.4]
  assign ridx_gray_io_d = _T_92 ^ _GEN_17; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310642.4]
  assign ridx_gray_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310643.4]
  assign AsyncValidSync_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310646.4]
  assign AsyncValidSync_reset = reset | _T_109; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310647.4 AsyncQueue.scala 157:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310657.4]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 160:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310662.4]
  assign AsyncValidSync_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310649.4]
  assign AsyncValidSync_1_reset = reset | _T_109; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310650.4 AsyncQueue.scala 158:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310661.4]
  assign AsyncValidSync_1_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 162:25:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310664.4]
  assign AsyncValidSync_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310652.4]
  assign AsyncValidSync_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310653.4]
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 163:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310665.4]
  assign AsyncResetRegVec_w1_i0_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310682.4]
  assign AsyncResetRegVec_w1_i0_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310683.4]
  assign AsyncResetRegVec_w1_i0_io_d = io_async_widx == io_async_ridx; // @[AsyncResetReg.scala 99:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310684.4]
  assign AsyncResetRegVec_w1_i0_io_en = 1'h1; // @[AsyncResetReg.scala 100:15:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310685.4]
endmodule
module AXI4AsyncCrossingSource( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310687.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310688.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310689.4]
  output        auto_in_aw_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_in_aw_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_in_aw_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [31:0] auto_in_aw_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_in_aw_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_in_w_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_in_w_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_in_w_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [7:0]  auto_in_w_bits_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_in_w_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_in_b_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_in_b_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_in_b_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_in_b_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_in_ar_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_in_ar_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_in_ar_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [31:0] auto_in_ar_bits_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_in_ar_bits_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_in_r_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_in_r_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_in_r_bits_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_in_r_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_in_r_bits_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_in_r_bits_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_aw_mem_0_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_aw_mem_0_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_0_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_aw_mem_0_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_mem_0_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_0_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_0_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_0_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_aw_mem_1_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_aw_mem_1_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_1_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_aw_mem_1_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_mem_1_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_1_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_1_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_1_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_aw_mem_2_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_aw_mem_2_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_2_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_aw_mem_2_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_mem_2_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_2_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_2_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_2_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_aw_mem_3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_aw_mem_3_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_3_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_aw_mem_3_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_mem_3_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_3_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_3_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_3_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_aw_mem_4_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_aw_mem_4_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_4_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_aw_mem_4_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_mem_4_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_4_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_4_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_4_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_aw_mem_5_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_aw_mem_5_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_5_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_aw_mem_5_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_mem_5_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_5_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_5_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_5_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_aw_mem_6_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_aw_mem_6_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_6_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_aw_mem_6_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_mem_6_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_6_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_6_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_6_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_aw_mem_7_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_aw_mem_7_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_7_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_aw_mem_7_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_mem_7_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_7_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_aw_mem_7_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_mem_7_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_aw_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_aw_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_aw_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_aw_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_aw_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_out_w_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_w_mem_0_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_out_w_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_w_mem_1_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_out_w_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_w_mem_2_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_out_w_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_w_mem_3_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_out_w_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_w_mem_4_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_out_w_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_w_mem_5_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_out_w_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_w_mem_6_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [63:0] auto_out_w_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_w_mem_7_strb, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_w_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_w_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_w_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_w_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_w_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_b_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_b_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_b_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_b_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_b_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_b_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_b_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_b_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_b_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_b_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_b_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_b_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_b_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_b_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_ar_mem_0_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_ar_mem_0_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_0_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_ar_mem_0_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_mem_0_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_0_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_0_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_0_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_ar_mem_1_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_ar_mem_1_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_1_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_ar_mem_1_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_mem_1_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_1_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_1_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_1_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_ar_mem_2_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_ar_mem_2_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_2_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_ar_mem_2_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_mem_2_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_2_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_2_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_2_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_ar_mem_3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_ar_mem_3_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_3_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_ar_mem_3_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_mem_3_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_3_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_3_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_3_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_ar_mem_4_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_ar_mem_4_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_4_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_ar_mem_4_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_mem_4_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_4_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_4_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_4_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_ar_mem_5_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_ar_mem_5_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_5_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_ar_mem_5_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_mem_5_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_5_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_5_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_5_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_ar_mem_6_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_ar_mem_6_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_6_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_ar_mem_6_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_mem_6_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_6_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_6_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_6_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [31:0] auto_out_ar_mem_7_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [7:0]  auto_out_ar_mem_7_len, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_7_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [1:0]  auto_out_ar_mem_7_burst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_mem_7_lock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_7_cache, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [2:0]  auto_out_ar_mem_7_prot, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_mem_7_qos, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_ar_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_ar_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_ar_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_ar_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_ar_safe_sink_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_mem_0_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_out_r_mem_0_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_r_mem_0_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_mem_0_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_mem_1_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_out_r_mem_1_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_r_mem_1_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_mem_1_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_mem_2_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_out_r_mem_2_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_r_mem_2_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_mem_2_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_mem_3_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_out_r_mem_3_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_r_mem_3_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_mem_3_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_mem_4_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_out_r_mem_4_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_r_mem_4_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_mem_4_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_mem_5_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_out_r_mem_5_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_r_mem_5_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_mem_5_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_mem_6_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_out_r_mem_6_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_r_mem_6_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_mem_6_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_mem_7_id, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [63:0] auto_out_r_mem_7_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [1:0]  auto_out_r_mem_7_resp, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_mem_7_last, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output [3:0]  auto_out_r_ridx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input  [3:0]  auto_out_r_widx, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_r_safe_ridx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_safe_widx_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  input         auto_out_r_safe_source_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
  output        auto_out_r_safe_sink_reset_n // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310690.4]
);
  wire  AsyncQueueSource_clock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_reset; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_enq_ready; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_enq_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_enq_bits_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_enq_bits_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_enq_bits_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_enq_bits_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_enq_bits_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_enq_bits_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_enq_bits_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_enq_bits_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_enq_bits_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_0_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_async_mem_0_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_async_mem_0_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_0_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_async_mem_0_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_mem_0_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_0_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_0_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_0_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_1_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_async_mem_1_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_async_mem_1_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_1_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_async_mem_1_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_mem_1_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_1_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_1_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_1_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_2_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_async_mem_2_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_async_mem_2_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_2_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_async_mem_2_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_mem_2_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_2_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_2_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_2_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_3_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_async_mem_3_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_async_mem_3_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_3_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_async_mem_3_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_mem_3_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_3_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_3_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_3_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_4_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_async_mem_4_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_async_mem_4_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_4_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_async_mem_4_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_mem_4_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_4_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_4_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_4_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_5_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_async_mem_5_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_async_mem_5_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_5_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_async_mem_5_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_mem_5_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_5_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_5_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_5_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_6_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_async_mem_6_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_async_mem_6_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_6_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_async_mem_6_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_mem_6_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_6_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_6_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_6_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_7_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [31:0] AsyncQueueSource_io_async_mem_7_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [7:0] AsyncQueueSource_io_async_mem_7_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_7_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [1:0] AsyncQueueSource_io_async_mem_7_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_mem_7_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_7_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [2:0] AsyncQueueSource_io_async_mem_7_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_mem_7_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_ridx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire [3:0] AsyncQueueSource_io_async_widx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_safe_ridx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_safe_widx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_safe_source_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
  wire  AsyncQueueSource_1_clock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_reset; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_enq_ready; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_enq_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_enq_bits_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_enq_bits_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_enq_bits_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_enq_bits_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_enq_bits_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_enq_bits_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_enq_bits_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_enq_bits_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_enq_bits_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_0_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_async_mem_0_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_async_mem_0_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_0_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_0_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_mem_0_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_0_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_0_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_0_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_1_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_async_mem_1_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_async_mem_1_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_1_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_1_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_mem_1_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_1_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_1_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_1_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_2_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_async_mem_2_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_async_mem_2_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_2_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_2_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_mem_2_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_2_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_2_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_2_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_3_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_async_mem_3_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_async_mem_3_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_3_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_3_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_mem_3_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_3_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_3_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_3_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_4_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_async_mem_4_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_async_mem_4_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_4_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_4_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_mem_4_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_4_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_4_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_4_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_5_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_async_mem_5_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_async_mem_5_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_5_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_5_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_mem_5_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_5_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_5_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_5_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_6_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_async_mem_6_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_async_mem_6_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_6_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_6_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_mem_6_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_6_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_6_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_6_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_7_id; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [31:0] AsyncQueueSource_1_io_async_mem_7_addr; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [7:0] AsyncQueueSource_1_io_async_mem_7_len; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_7_size; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [1:0] AsyncQueueSource_1_io_async_mem_7_burst; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_mem_7_lock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_7_cache; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [2:0] AsyncQueueSource_1_io_async_mem_7_prot; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_mem_7_qos; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_ridx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire [3:0] AsyncQueueSource_1_io_async_widx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_safe_ridx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_safe_widx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_safe_source_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_1_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
  wire  AsyncQueueSource_2_clock; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_reset; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_enq_ready; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_enq_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_enq_bits_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_enq_bits_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_enq_bits_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_async_mem_0_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_async_mem_0_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_mem_0_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_async_mem_1_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_async_mem_1_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_mem_1_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_async_mem_2_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_async_mem_2_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_mem_2_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_async_mem_3_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_async_mem_3_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_mem_3_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_async_mem_4_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_async_mem_4_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_mem_4_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_async_mem_5_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_async_mem_5_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_mem_5_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_async_mem_6_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_async_mem_6_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_mem_6_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [63:0] AsyncQueueSource_2_io_async_mem_7_data; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [7:0] AsyncQueueSource_2_io_async_mem_7_strb; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_mem_7_last; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [3:0] AsyncQueueSource_2_io_async_ridx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire [3:0] AsyncQueueSource_2_io_async_widx; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_safe_ridx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_safe_widx_valid; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_safe_source_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSource_2_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
  wire  AsyncQueueSink_clock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_reset; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_deq_ready; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_deq_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_deq_bits_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_deq_bits_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_deq_bits_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_deq_bits_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_mem_0_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_async_mem_0_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_async_mem_0_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_mem_0_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_mem_1_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_async_mem_1_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_async_mem_1_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_mem_1_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_mem_2_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_async_mem_2_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_async_mem_2_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_mem_2_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_mem_3_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_async_mem_3_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_async_mem_3_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_mem_3_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_mem_4_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_async_mem_4_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_async_mem_4_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_mem_4_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_mem_5_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_async_mem_5_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_async_mem_5_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_mem_5_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_mem_6_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_async_mem_6_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_async_mem_6_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_mem_6_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_mem_7_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [63:0] AsyncQueueSink_io_async_mem_7_data; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [1:0] AsyncQueueSink_io_async_mem_7_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_mem_7_last; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_ridx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire [3:0] AsyncQueueSink_io_async_widx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_safe_widx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
  wire  AsyncQueueSink_1_clock; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire  AsyncQueueSink_1_reset; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire  AsyncQueueSink_1_io_deq_ready; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire  AsyncQueueSink_1_io_deq_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_deq_bits_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_deq_bits_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_0_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_0_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_1_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_1_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_2_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_2_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_3_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_3_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_4_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_4_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_5_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_5_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_6_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_6_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_mem_7_id; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [1:0] AsyncQueueSink_1_io_async_mem_7_resp; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_ridx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire [3:0] AsyncQueueSink_1_io_async_widx; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire  AsyncQueueSink_1_io_async_safe_ridx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire  AsyncQueueSink_1_io_async_safe_widx_valid; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire  AsyncQueueSink_1_io_async_safe_source_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  wire  AsyncQueueSink_1_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
  AsyncQueueSource_5 AsyncQueueSource ( // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310701.4]
    .clock(AsyncQueueSource_clock),
    .reset(AsyncQueueSource_reset),
    .io_enq_ready(AsyncQueueSource_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_io_enq_valid),
    .io_enq_bits_id(AsyncQueueSource_io_enq_bits_id),
    .io_enq_bits_addr(AsyncQueueSource_io_enq_bits_addr),
    .io_enq_bits_len(AsyncQueueSource_io_enq_bits_len),
    .io_enq_bits_size(AsyncQueueSource_io_enq_bits_size),
    .io_enq_bits_burst(AsyncQueueSource_io_enq_bits_burst),
    .io_enq_bits_lock(AsyncQueueSource_io_enq_bits_lock),
    .io_enq_bits_cache(AsyncQueueSource_io_enq_bits_cache),
    .io_enq_bits_prot(AsyncQueueSource_io_enq_bits_prot),
    .io_enq_bits_qos(AsyncQueueSource_io_enq_bits_qos),
    .io_async_mem_0_id(AsyncQueueSource_io_async_mem_0_id),
    .io_async_mem_0_addr(AsyncQueueSource_io_async_mem_0_addr),
    .io_async_mem_0_len(AsyncQueueSource_io_async_mem_0_len),
    .io_async_mem_0_size(AsyncQueueSource_io_async_mem_0_size),
    .io_async_mem_0_burst(AsyncQueueSource_io_async_mem_0_burst),
    .io_async_mem_0_lock(AsyncQueueSource_io_async_mem_0_lock),
    .io_async_mem_0_cache(AsyncQueueSource_io_async_mem_0_cache),
    .io_async_mem_0_prot(AsyncQueueSource_io_async_mem_0_prot),
    .io_async_mem_0_qos(AsyncQueueSource_io_async_mem_0_qos),
    .io_async_mem_1_id(AsyncQueueSource_io_async_mem_1_id),
    .io_async_mem_1_addr(AsyncQueueSource_io_async_mem_1_addr),
    .io_async_mem_1_len(AsyncQueueSource_io_async_mem_1_len),
    .io_async_mem_1_size(AsyncQueueSource_io_async_mem_1_size),
    .io_async_mem_1_burst(AsyncQueueSource_io_async_mem_1_burst),
    .io_async_mem_1_lock(AsyncQueueSource_io_async_mem_1_lock),
    .io_async_mem_1_cache(AsyncQueueSource_io_async_mem_1_cache),
    .io_async_mem_1_prot(AsyncQueueSource_io_async_mem_1_prot),
    .io_async_mem_1_qos(AsyncQueueSource_io_async_mem_1_qos),
    .io_async_mem_2_id(AsyncQueueSource_io_async_mem_2_id),
    .io_async_mem_2_addr(AsyncQueueSource_io_async_mem_2_addr),
    .io_async_mem_2_len(AsyncQueueSource_io_async_mem_2_len),
    .io_async_mem_2_size(AsyncQueueSource_io_async_mem_2_size),
    .io_async_mem_2_burst(AsyncQueueSource_io_async_mem_2_burst),
    .io_async_mem_2_lock(AsyncQueueSource_io_async_mem_2_lock),
    .io_async_mem_2_cache(AsyncQueueSource_io_async_mem_2_cache),
    .io_async_mem_2_prot(AsyncQueueSource_io_async_mem_2_prot),
    .io_async_mem_2_qos(AsyncQueueSource_io_async_mem_2_qos),
    .io_async_mem_3_id(AsyncQueueSource_io_async_mem_3_id),
    .io_async_mem_3_addr(AsyncQueueSource_io_async_mem_3_addr),
    .io_async_mem_3_len(AsyncQueueSource_io_async_mem_3_len),
    .io_async_mem_3_size(AsyncQueueSource_io_async_mem_3_size),
    .io_async_mem_3_burst(AsyncQueueSource_io_async_mem_3_burst),
    .io_async_mem_3_lock(AsyncQueueSource_io_async_mem_3_lock),
    .io_async_mem_3_cache(AsyncQueueSource_io_async_mem_3_cache),
    .io_async_mem_3_prot(AsyncQueueSource_io_async_mem_3_prot),
    .io_async_mem_3_qos(AsyncQueueSource_io_async_mem_3_qos),
    .io_async_mem_4_id(AsyncQueueSource_io_async_mem_4_id),
    .io_async_mem_4_addr(AsyncQueueSource_io_async_mem_4_addr),
    .io_async_mem_4_len(AsyncQueueSource_io_async_mem_4_len),
    .io_async_mem_4_size(AsyncQueueSource_io_async_mem_4_size),
    .io_async_mem_4_burst(AsyncQueueSource_io_async_mem_4_burst),
    .io_async_mem_4_lock(AsyncQueueSource_io_async_mem_4_lock),
    .io_async_mem_4_cache(AsyncQueueSource_io_async_mem_4_cache),
    .io_async_mem_4_prot(AsyncQueueSource_io_async_mem_4_prot),
    .io_async_mem_4_qos(AsyncQueueSource_io_async_mem_4_qos),
    .io_async_mem_5_id(AsyncQueueSource_io_async_mem_5_id),
    .io_async_mem_5_addr(AsyncQueueSource_io_async_mem_5_addr),
    .io_async_mem_5_len(AsyncQueueSource_io_async_mem_5_len),
    .io_async_mem_5_size(AsyncQueueSource_io_async_mem_5_size),
    .io_async_mem_5_burst(AsyncQueueSource_io_async_mem_5_burst),
    .io_async_mem_5_lock(AsyncQueueSource_io_async_mem_5_lock),
    .io_async_mem_5_cache(AsyncQueueSource_io_async_mem_5_cache),
    .io_async_mem_5_prot(AsyncQueueSource_io_async_mem_5_prot),
    .io_async_mem_5_qos(AsyncQueueSource_io_async_mem_5_qos),
    .io_async_mem_6_id(AsyncQueueSource_io_async_mem_6_id),
    .io_async_mem_6_addr(AsyncQueueSource_io_async_mem_6_addr),
    .io_async_mem_6_len(AsyncQueueSource_io_async_mem_6_len),
    .io_async_mem_6_size(AsyncQueueSource_io_async_mem_6_size),
    .io_async_mem_6_burst(AsyncQueueSource_io_async_mem_6_burst),
    .io_async_mem_6_lock(AsyncQueueSource_io_async_mem_6_lock),
    .io_async_mem_6_cache(AsyncQueueSource_io_async_mem_6_cache),
    .io_async_mem_6_prot(AsyncQueueSource_io_async_mem_6_prot),
    .io_async_mem_6_qos(AsyncQueueSource_io_async_mem_6_qos),
    .io_async_mem_7_id(AsyncQueueSource_io_async_mem_7_id),
    .io_async_mem_7_addr(AsyncQueueSource_io_async_mem_7_addr),
    .io_async_mem_7_len(AsyncQueueSource_io_async_mem_7_len),
    .io_async_mem_7_size(AsyncQueueSource_io_async_mem_7_size),
    .io_async_mem_7_burst(AsyncQueueSource_io_async_mem_7_burst),
    .io_async_mem_7_lock(AsyncQueueSource_io_async_mem_7_lock),
    .io_async_mem_7_cache(AsyncQueueSource_io_async_mem_7_cache),
    .io_async_mem_7_prot(AsyncQueueSource_io_async_mem_7_prot),
    .io_async_mem_7_qos(AsyncQueueSource_io_async_mem_7_qos),
    .io_async_ridx(AsyncQueueSource_io_async_ridx),
    .io_async_widx(AsyncQueueSource_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource_5 AsyncQueueSource_1 ( // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310708.4]
    .clock(AsyncQueueSource_1_clock),
    .reset(AsyncQueueSource_1_reset),
    .io_enq_ready(AsyncQueueSource_1_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_1_io_enq_valid),
    .io_enq_bits_id(AsyncQueueSource_1_io_enq_bits_id),
    .io_enq_bits_addr(AsyncQueueSource_1_io_enq_bits_addr),
    .io_enq_bits_len(AsyncQueueSource_1_io_enq_bits_len),
    .io_enq_bits_size(AsyncQueueSource_1_io_enq_bits_size),
    .io_enq_bits_burst(AsyncQueueSource_1_io_enq_bits_burst),
    .io_enq_bits_lock(AsyncQueueSource_1_io_enq_bits_lock),
    .io_enq_bits_cache(AsyncQueueSource_1_io_enq_bits_cache),
    .io_enq_bits_prot(AsyncQueueSource_1_io_enq_bits_prot),
    .io_enq_bits_qos(AsyncQueueSource_1_io_enq_bits_qos),
    .io_async_mem_0_id(AsyncQueueSource_1_io_async_mem_0_id),
    .io_async_mem_0_addr(AsyncQueueSource_1_io_async_mem_0_addr),
    .io_async_mem_0_len(AsyncQueueSource_1_io_async_mem_0_len),
    .io_async_mem_0_size(AsyncQueueSource_1_io_async_mem_0_size),
    .io_async_mem_0_burst(AsyncQueueSource_1_io_async_mem_0_burst),
    .io_async_mem_0_lock(AsyncQueueSource_1_io_async_mem_0_lock),
    .io_async_mem_0_cache(AsyncQueueSource_1_io_async_mem_0_cache),
    .io_async_mem_0_prot(AsyncQueueSource_1_io_async_mem_0_prot),
    .io_async_mem_0_qos(AsyncQueueSource_1_io_async_mem_0_qos),
    .io_async_mem_1_id(AsyncQueueSource_1_io_async_mem_1_id),
    .io_async_mem_1_addr(AsyncQueueSource_1_io_async_mem_1_addr),
    .io_async_mem_1_len(AsyncQueueSource_1_io_async_mem_1_len),
    .io_async_mem_1_size(AsyncQueueSource_1_io_async_mem_1_size),
    .io_async_mem_1_burst(AsyncQueueSource_1_io_async_mem_1_burst),
    .io_async_mem_1_lock(AsyncQueueSource_1_io_async_mem_1_lock),
    .io_async_mem_1_cache(AsyncQueueSource_1_io_async_mem_1_cache),
    .io_async_mem_1_prot(AsyncQueueSource_1_io_async_mem_1_prot),
    .io_async_mem_1_qos(AsyncQueueSource_1_io_async_mem_1_qos),
    .io_async_mem_2_id(AsyncQueueSource_1_io_async_mem_2_id),
    .io_async_mem_2_addr(AsyncQueueSource_1_io_async_mem_2_addr),
    .io_async_mem_2_len(AsyncQueueSource_1_io_async_mem_2_len),
    .io_async_mem_2_size(AsyncQueueSource_1_io_async_mem_2_size),
    .io_async_mem_2_burst(AsyncQueueSource_1_io_async_mem_2_burst),
    .io_async_mem_2_lock(AsyncQueueSource_1_io_async_mem_2_lock),
    .io_async_mem_2_cache(AsyncQueueSource_1_io_async_mem_2_cache),
    .io_async_mem_2_prot(AsyncQueueSource_1_io_async_mem_2_prot),
    .io_async_mem_2_qos(AsyncQueueSource_1_io_async_mem_2_qos),
    .io_async_mem_3_id(AsyncQueueSource_1_io_async_mem_3_id),
    .io_async_mem_3_addr(AsyncQueueSource_1_io_async_mem_3_addr),
    .io_async_mem_3_len(AsyncQueueSource_1_io_async_mem_3_len),
    .io_async_mem_3_size(AsyncQueueSource_1_io_async_mem_3_size),
    .io_async_mem_3_burst(AsyncQueueSource_1_io_async_mem_3_burst),
    .io_async_mem_3_lock(AsyncQueueSource_1_io_async_mem_3_lock),
    .io_async_mem_3_cache(AsyncQueueSource_1_io_async_mem_3_cache),
    .io_async_mem_3_prot(AsyncQueueSource_1_io_async_mem_3_prot),
    .io_async_mem_3_qos(AsyncQueueSource_1_io_async_mem_3_qos),
    .io_async_mem_4_id(AsyncQueueSource_1_io_async_mem_4_id),
    .io_async_mem_4_addr(AsyncQueueSource_1_io_async_mem_4_addr),
    .io_async_mem_4_len(AsyncQueueSource_1_io_async_mem_4_len),
    .io_async_mem_4_size(AsyncQueueSource_1_io_async_mem_4_size),
    .io_async_mem_4_burst(AsyncQueueSource_1_io_async_mem_4_burst),
    .io_async_mem_4_lock(AsyncQueueSource_1_io_async_mem_4_lock),
    .io_async_mem_4_cache(AsyncQueueSource_1_io_async_mem_4_cache),
    .io_async_mem_4_prot(AsyncQueueSource_1_io_async_mem_4_prot),
    .io_async_mem_4_qos(AsyncQueueSource_1_io_async_mem_4_qos),
    .io_async_mem_5_id(AsyncQueueSource_1_io_async_mem_5_id),
    .io_async_mem_5_addr(AsyncQueueSource_1_io_async_mem_5_addr),
    .io_async_mem_5_len(AsyncQueueSource_1_io_async_mem_5_len),
    .io_async_mem_5_size(AsyncQueueSource_1_io_async_mem_5_size),
    .io_async_mem_5_burst(AsyncQueueSource_1_io_async_mem_5_burst),
    .io_async_mem_5_lock(AsyncQueueSource_1_io_async_mem_5_lock),
    .io_async_mem_5_cache(AsyncQueueSource_1_io_async_mem_5_cache),
    .io_async_mem_5_prot(AsyncQueueSource_1_io_async_mem_5_prot),
    .io_async_mem_5_qos(AsyncQueueSource_1_io_async_mem_5_qos),
    .io_async_mem_6_id(AsyncQueueSource_1_io_async_mem_6_id),
    .io_async_mem_6_addr(AsyncQueueSource_1_io_async_mem_6_addr),
    .io_async_mem_6_len(AsyncQueueSource_1_io_async_mem_6_len),
    .io_async_mem_6_size(AsyncQueueSource_1_io_async_mem_6_size),
    .io_async_mem_6_burst(AsyncQueueSource_1_io_async_mem_6_burst),
    .io_async_mem_6_lock(AsyncQueueSource_1_io_async_mem_6_lock),
    .io_async_mem_6_cache(AsyncQueueSource_1_io_async_mem_6_cache),
    .io_async_mem_6_prot(AsyncQueueSource_1_io_async_mem_6_prot),
    .io_async_mem_6_qos(AsyncQueueSource_1_io_async_mem_6_qos),
    .io_async_mem_7_id(AsyncQueueSource_1_io_async_mem_7_id),
    .io_async_mem_7_addr(AsyncQueueSource_1_io_async_mem_7_addr),
    .io_async_mem_7_len(AsyncQueueSource_1_io_async_mem_7_len),
    .io_async_mem_7_size(AsyncQueueSource_1_io_async_mem_7_size),
    .io_async_mem_7_burst(AsyncQueueSource_1_io_async_mem_7_burst),
    .io_async_mem_7_lock(AsyncQueueSource_1_io_async_mem_7_lock),
    .io_async_mem_7_cache(AsyncQueueSource_1_io_async_mem_7_cache),
    .io_async_mem_7_prot(AsyncQueueSource_1_io_async_mem_7_prot),
    .io_async_mem_7_qos(AsyncQueueSource_1_io_async_mem_7_qos),
    .io_async_ridx(AsyncQueueSource_1_io_async_ridx),
    .io_async_widx(AsyncQueueSource_1_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_1_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_1_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_1_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_1_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource_7 AsyncQueueSource_2 ( // @[AsyncQueue.scala 192:24:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310715.4]
    .clock(AsyncQueueSource_2_clock),
    .reset(AsyncQueueSource_2_reset),
    .io_enq_ready(AsyncQueueSource_2_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_2_io_enq_valid),
    .io_enq_bits_data(AsyncQueueSource_2_io_enq_bits_data),
    .io_enq_bits_strb(AsyncQueueSource_2_io_enq_bits_strb),
    .io_enq_bits_last(AsyncQueueSource_2_io_enq_bits_last),
    .io_async_mem_0_data(AsyncQueueSource_2_io_async_mem_0_data),
    .io_async_mem_0_strb(AsyncQueueSource_2_io_async_mem_0_strb),
    .io_async_mem_0_last(AsyncQueueSource_2_io_async_mem_0_last),
    .io_async_mem_1_data(AsyncQueueSource_2_io_async_mem_1_data),
    .io_async_mem_1_strb(AsyncQueueSource_2_io_async_mem_1_strb),
    .io_async_mem_1_last(AsyncQueueSource_2_io_async_mem_1_last),
    .io_async_mem_2_data(AsyncQueueSource_2_io_async_mem_2_data),
    .io_async_mem_2_strb(AsyncQueueSource_2_io_async_mem_2_strb),
    .io_async_mem_2_last(AsyncQueueSource_2_io_async_mem_2_last),
    .io_async_mem_3_data(AsyncQueueSource_2_io_async_mem_3_data),
    .io_async_mem_3_strb(AsyncQueueSource_2_io_async_mem_3_strb),
    .io_async_mem_3_last(AsyncQueueSource_2_io_async_mem_3_last),
    .io_async_mem_4_data(AsyncQueueSource_2_io_async_mem_4_data),
    .io_async_mem_4_strb(AsyncQueueSource_2_io_async_mem_4_strb),
    .io_async_mem_4_last(AsyncQueueSource_2_io_async_mem_4_last),
    .io_async_mem_5_data(AsyncQueueSource_2_io_async_mem_5_data),
    .io_async_mem_5_strb(AsyncQueueSource_2_io_async_mem_5_strb),
    .io_async_mem_5_last(AsyncQueueSource_2_io_async_mem_5_last),
    .io_async_mem_6_data(AsyncQueueSource_2_io_async_mem_6_data),
    .io_async_mem_6_strb(AsyncQueueSource_2_io_async_mem_6_strb),
    .io_async_mem_6_last(AsyncQueueSource_2_io_async_mem_6_last),
    .io_async_mem_7_data(AsyncQueueSource_2_io_async_mem_7_data),
    .io_async_mem_7_strb(AsyncQueueSource_2_io_async_mem_7_strb),
    .io_async_mem_7_last(AsyncQueueSource_2_io_async_mem_7_last),
    .io_async_ridx(AsyncQueueSource_2_io_async_ridx),
    .io_async_widx(AsyncQueueSource_2_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_2_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_2_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_2_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_2_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink_6 AsyncQueueSink ( // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310722.4]
    .clock(AsyncQueueSink_clock),
    .reset(AsyncQueueSink_reset),
    .io_deq_ready(AsyncQueueSink_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_io_deq_valid),
    .io_deq_bits_id(AsyncQueueSink_io_deq_bits_id),
    .io_deq_bits_data(AsyncQueueSink_io_deq_bits_data),
    .io_deq_bits_resp(AsyncQueueSink_io_deq_bits_resp),
    .io_deq_bits_last(AsyncQueueSink_io_deq_bits_last),
    .io_async_mem_0_id(AsyncQueueSink_io_async_mem_0_id),
    .io_async_mem_0_data(AsyncQueueSink_io_async_mem_0_data),
    .io_async_mem_0_resp(AsyncQueueSink_io_async_mem_0_resp),
    .io_async_mem_0_last(AsyncQueueSink_io_async_mem_0_last),
    .io_async_mem_1_id(AsyncQueueSink_io_async_mem_1_id),
    .io_async_mem_1_data(AsyncQueueSink_io_async_mem_1_data),
    .io_async_mem_1_resp(AsyncQueueSink_io_async_mem_1_resp),
    .io_async_mem_1_last(AsyncQueueSink_io_async_mem_1_last),
    .io_async_mem_2_id(AsyncQueueSink_io_async_mem_2_id),
    .io_async_mem_2_data(AsyncQueueSink_io_async_mem_2_data),
    .io_async_mem_2_resp(AsyncQueueSink_io_async_mem_2_resp),
    .io_async_mem_2_last(AsyncQueueSink_io_async_mem_2_last),
    .io_async_mem_3_id(AsyncQueueSink_io_async_mem_3_id),
    .io_async_mem_3_data(AsyncQueueSink_io_async_mem_3_data),
    .io_async_mem_3_resp(AsyncQueueSink_io_async_mem_3_resp),
    .io_async_mem_3_last(AsyncQueueSink_io_async_mem_3_last),
    .io_async_mem_4_id(AsyncQueueSink_io_async_mem_4_id),
    .io_async_mem_4_data(AsyncQueueSink_io_async_mem_4_data),
    .io_async_mem_4_resp(AsyncQueueSink_io_async_mem_4_resp),
    .io_async_mem_4_last(AsyncQueueSink_io_async_mem_4_last),
    .io_async_mem_5_id(AsyncQueueSink_io_async_mem_5_id),
    .io_async_mem_5_data(AsyncQueueSink_io_async_mem_5_data),
    .io_async_mem_5_resp(AsyncQueueSink_io_async_mem_5_resp),
    .io_async_mem_5_last(AsyncQueueSink_io_async_mem_5_last),
    .io_async_mem_6_id(AsyncQueueSink_io_async_mem_6_id),
    .io_async_mem_6_data(AsyncQueueSink_io_async_mem_6_data),
    .io_async_mem_6_resp(AsyncQueueSink_io_async_mem_6_resp),
    .io_async_mem_6_last(AsyncQueueSink_io_async_mem_6_last),
    .io_async_mem_7_id(AsyncQueueSink_io_async_mem_7_id),
    .io_async_mem_7_data(AsyncQueueSink_io_async_mem_7_data),
    .io_async_mem_7_resp(AsyncQueueSink_io_async_mem_7_resp),
    .io_async_mem_7_last(AsyncQueueSink_io_async_mem_7_last),
    .io_async_ridx(AsyncQueueSink_io_async_ridx),
    .io_async_widx(AsyncQueueSink_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink_7 AsyncQueueSink_1 ( // @[AsyncQueue.scala 183:22:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310740.4]
    .clock(AsyncQueueSink_1_clock),
    .reset(AsyncQueueSink_1_reset),
    .io_deq_ready(AsyncQueueSink_1_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_1_io_deq_valid),
    .io_deq_bits_id(AsyncQueueSink_1_io_deq_bits_id),
    .io_deq_bits_resp(AsyncQueueSink_1_io_deq_bits_resp),
    .io_async_mem_0_id(AsyncQueueSink_1_io_async_mem_0_id),
    .io_async_mem_0_resp(AsyncQueueSink_1_io_async_mem_0_resp),
    .io_async_mem_1_id(AsyncQueueSink_1_io_async_mem_1_id),
    .io_async_mem_1_resp(AsyncQueueSink_1_io_async_mem_1_resp),
    .io_async_mem_2_id(AsyncQueueSink_1_io_async_mem_2_id),
    .io_async_mem_2_resp(AsyncQueueSink_1_io_async_mem_2_resp),
    .io_async_mem_3_id(AsyncQueueSink_1_io_async_mem_3_id),
    .io_async_mem_3_resp(AsyncQueueSink_1_io_async_mem_3_resp),
    .io_async_mem_4_id(AsyncQueueSink_1_io_async_mem_4_id),
    .io_async_mem_4_resp(AsyncQueueSink_1_io_async_mem_4_resp),
    .io_async_mem_5_id(AsyncQueueSink_1_io_async_mem_5_id),
    .io_async_mem_5_resp(AsyncQueueSink_1_io_async_mem_5_resp),
    .io_async_mem_6_id(AsyncQueueSink_1_io_async_mem_6_id),
    .io_async_mem_6_resp(AsyncQueueSink_1_io_async_mem_6_resp),
    .io_async_mem_7_id(AsyncQueueSink_1_io_async_mem_7_id),
    .io_async_mem_7_resp(AsyncQueueSink_1_io_async_mem_7_resp),
    .io_async_ridx(AsyncQueueSink_1_io_async_ridx),
    .io_async_widx(AsyncQueueSink_1_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_1_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_1_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_1_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_1_io_async_safe_sink_reset_n)
  );
  assign auto_in_aw_ready = AsyncQueueSource_1_io_enq_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_w_ready = AsyncQueueSource_2_io_enq_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_b_valid = AsyncQueueSink_1_io_deq_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_b_bits_id = AsyncQueueSink_1_io_deq_bits_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_b_bits_resp = AsyncQueueSink_1_io_deq_bits_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_ar_ready = AsyncQueueSource_io_enq_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_r_valid = AsyncQueueSink_io_deq_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_r_bits_id = AsyncQueueSink_io_deq_bits_id; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_r_bits_data = AsyncQueueSink_io_deq_bits_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_r_bits_resp = AsyncQueueSink_io_deq_bits_resp; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_in_r_bits_last = AsyncQueueSink_io_deq_bits_last; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310700.4]
  assign auto_out_aw_mem_0_id = AsyncQueueSource_1_io_async_mem_0_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_0_addr = AsyncQueueSource_1_io_async_mem_0_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_0_len = AsyncQueueSource_1_io_async_mem_0_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_0_size = AsyncQueueSource_1_io_async_mem_0_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_0_burst = AsyncQueueSource_1_io_async_mem_0_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_0_lock = AsyncQueueSource_1_io_async_mem_0_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_0_cache = AsyncQueueSource_1_io_async_mem_0_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_0_prot = AsyncQueueSource_1_io_async_mem_0_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_0_qos = AsyncQueueSource_1_io_async_mem_0_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_id = AsyncQueueSource_1_io_async_mem_1_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_addr = AsyncQueueSource_1_io_async_mem_1_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_len = AsyncQueueSource_1_io_async_mem_1_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_size = AsyncQueueSource_1_io_async_mem_1_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_burst = AsyncQueueSource_1_io_async_mem_1_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_lock = AsyncQueueSource_1_io_async_mem_1_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_cache = AsyncQueueSource_1_io_async_mem_1_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_prot = AsyncQueueSource_1_io_async_mem_1_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_1_qos = AsyncQueueSource_1_io_async_mem_1_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_id = AsyncQueueSource_1_io_async_mem_2_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_addr = AsyncQueueSource_1_io_async_mem_2_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_len = AsyncQueueSource_1_io_async_mem_2_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_size = AsyncQueueSource_1_io_async_mem_2_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_burst = AsyncQueueSource_1_io_async_mem_2_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_lock = AsyncQueueSource_1_io_async_mem_2_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_cache = AsyncQueueSource_1_io_async_mem_2_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_prot = AsyncQueueSource_1_io_async_mem_2_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_2_qos = AsyncQueueSource_1_io_async_mem_2_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_id = AsyncQueueSource_1_io_async_mem_3_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_addr = AsyncQueueSource_1_io_async_mem_3_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_len = AsyncQueueSource_1_io_async_mem_3_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_size = AsyncQueueSource_1_io_async_mem_3_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_burst = AsyncQueueSource_1_io_async_mem_3_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_lock = AsyncQueueSource_1_io_async_mem_3_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_cache = AsyncQueueSource_1_io_async_mem_3_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_prot = AsyncQueueSource_1_io_async_mem_3_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_3_qos = AsyncQueueSource_1_io_async_mem_3_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_id = AsyncQueueSource_1_io_async_mem_4_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_addr = AsyncQueueSource_1_io_async_mem_4_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_len = AsyncQueueSource_1_io_async_mem_4_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_size = AsyncQueueSource_1_io_async_mem_4_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_burst = AsyncQueueSource_1_io_async_mem_4_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_lock = AsyncQueueSource_1_io_async_mem_4_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_cache = AsyncQueueSource_1_io_async_mem_4_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_prot = AsyncQueueSource_1_io_async_mem_4_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_4_qos = AsyncQueueSource_1_io_async_mem_4_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_id = AsyncQueueSource_1_io_async_mem_5_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_addr = AsyncQueueSource_1_io_async_mem_5_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_len = AsyncQueueSource_1_io_async_mem_5_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_size = AsyncQueueSource_1_io_async_mem_5_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_burst = AsyncQueueSource_1_io_async_mem_5_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_lock = AsyncQueueSource_1_io_async_mem_5_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_cache = AsyncQueueSource_1_io_async_mem_5_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_prot = AsyncQueueSource_1_io_async_mem_5_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_5_qos = AsyncQueueSource_1_io_async_mem_5_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_id = AsyncQueueSource_1_io_async_mem_6_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_addr = AsyncQueueSource_1_io_async_mem_6_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_len = AsyncQueueSource_1_io_async_mem_6_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_size = AsyncQueueSource_1_io_async_mem_6_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_burst = AsyncQueueSource_1_io_async_mem_6_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_lock = AsyncQueueSource_1_io_async_mem_6_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_cache = AsyncQueueSource_1_io_async_mem_6_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_prot = AsyncQueueSource_1_io_async_mem_6_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_6_qos = AsyncQueueSource_1_io_async_mem_6_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_id = AsyncQueueSource_1_io_async_mem_7_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_addr = AsyncQueueSource_1_io_async_mem_7_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_len = AsyncQueueSource_1_io_async_mem_7_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_size = AsyncQueueSource_1_io_async_mem_7_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_burst = AsyncQueueSource_1_io_async_mem_7_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_lock = AsyncQueueSource_1_io_async_mem_7_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_cache = AsyncQueueSource_1_io_async_mem_7_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_prot = AsyncQueueSource_1_io_async_mem_7_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_mem_7_qos = AsyncQueueSource_1_io_async_mem_7_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_widx = AsyncQueueSource_1_io_async_widx; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_safe_widx_valid = AsyncQueueSource_1_io_async_safe_widx_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_aw_safe_source_reset_n = AsyncQueueSource_1_io_async_safe_source_reset_n; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_0_data = AsyncQueueSource_2_io_async_mem_0_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_0_strb = AsyncQueueSource_2_io_async_mem_0_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_0_last = AsyncQueueSource_2_io_async_mem_0_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_1_data = AsyncQueueSource_2_io_async_mem_1_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_1_strb = AsyncQueueSource_2_io_async_mem_1_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_1_last = AsyncQueueSource_2_io_async_mem_1_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_2_data = AsyncQueueSource_2_io_async_mem_2_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_2_strb = AsyncQueueSource_2_io_async_mem_2_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_2_last = AsyncQueueSource_2_io_async_mem_2_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_3_data = AsyncQueueSource_2_io_async_mem_3_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_3_strb = AsyncQueueSource_2_io_async_mem_3_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_3_last = AsyncQueueSource_2_io_async_mem_3_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_4_data = AsyncQueueSource_2_io_async_mem_4_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_4_strb = AsyncQueueSource_2_io_async_mem_4_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_4_last = AsyncQueueSource_2_io_async_mem_4_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_5_data = AsyncQueueSource_2_io_async_mem_5_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_5_strb = AsyncQueueSource_2_io_async_mem_5_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_5_last = AsyncQueueSource_2_io_async_mem_5_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_6_data = AsyncQueueSource_2_io_async_mem_6_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_6_strb = AsyncQueueSource_2_io_async_mem_6_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_6_last = AsyncQueueSource_2_io_async_mem_6_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_7_data = AsyncQueueSource_2_io_async_mem_7_data; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_7_strb = AsyncQueueSource_2_io_async_mem_7_strb; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_mem_7_last = AsyncQueueSource_2_io_async_mem_7_last; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_widx = AsyncQueueSource_2_io_async_widx; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_safe_widx_valid = AsyncQueueSource_2_io_async_safe_widx_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_w_safe_source_reset_n = AsyncQueueSource_2_io_async_safe_source_reset_n; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_b_ridx = AsyncQueueSink_1_io_async_ridx; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_b_safe_ridx_valid = AsyncQueueSink_1_io_async_safe_ridx_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_b_safe_sink_reset_n = AsyncQueueSink_1_io_async_safe_sink_reset_n; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_id = AsyncQueueSource_io_async_mem_0_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_addr = AsyncQueueSource_io_async_mem_0_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_len = AsyncQueueSource_io_async_mem_0_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_size = AsyncQueueSource_io_async_mem_0_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_burst = AsyncQueueSource_io_async_mem_0_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_lock = AsyncQueueSource_io_async_mem_0_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_cache = AsyncQueueSource_io_async_mem_0_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_prot = AsyncQueueSource_io_async_mem_0_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_0_qos = AsyncQueueSource_io_async_mem_0_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_id = AsyncQueueSource_io_async_mem_1_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_addr = AsyncQueueSource_io_async_mem_1_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_len = AsyncQueueSource_io_async_mem_1_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_size = AsyncQueueSource_io_async_mem_1_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_burst = AsyncQueueSource_io_async_mem_1_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_lock = AsyncQueueSource_io_async_mem_1_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_cache = AsyncQueueSource_io_async_mem_1_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_prot = AsyncQueueSource_io_async_mem_1_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_1_qos = AsyncQueueSource_io_async_mem_1_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_id = AsyncQueueSource_io_async_mem_2_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_addr = AsyncQueueSource_io_async_mem_2_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_len = AsyncQueueSource_io_async_mem_2_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_size = AsyncQueueSource_io_async_mem_2_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_burst = AsyncQueueSource_io_async_mem_2_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_lock = AsyncQueueSource_io_async_mem_2_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_cache = AsyncQueueSource_io_async_mem_2_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_prot = AsyncQueueSource_io_async_mem_2_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_2_qos = AsyncQueueSource_io_async_mem_2_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_id = AsyncQueueSource_io_async_mem_3_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_addr = AsyncQueueSource_io_async_mem_3_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_len = AsyncQueueSource_io_async_mem_3_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_size = AsyncQueueSource_io_async_mem_3_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_burst = AsyncQueueSource_io_async_mem_3_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_lock = AsyncQueueSource_io_async_mem_3_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_cache = AsyncQueueSource_io_async_mem_3_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_prot = AsyncQueueSource_io_async_mem_3_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_3_qos = AsyncQueueSource_io_async_mem_3_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_id = AsyncQueueSource_io_async_mem_4_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_addr = AsyncQueueSource_io_async_mem_4_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_len = AsyncQueueSource_io_async_mem_4_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_size = AsyncQueueSource_io_async_mem_4_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_burst = AsyncQueueSource_io_async_mem_4_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_lock = AsyncQueueSource_io_async_mem_4_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_cache = AsyncQueueSource_io_async_mem_4_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_prot = AsyncQueueSource_io_async_mem_4_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_4_qos = AsyncQueueSource_io_async_mem_4_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_id = AsyncQueueSource_io_async_mem_5_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_addr = AsyncQueueSource_io_async_mem_5_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_len = AsyncQueueSource_io_async_mem_5_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_size = AsyncQueueSource_io_async_mem_5_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_burst = AsyncQueueSource_io_async_mem_5_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_lock = AsyncQueueSource_io_async_mem_5_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_cache = AsyncQueueSource_io_async_mem_5_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_prot = AsyncQueueSource_io_async_mem_5_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_5_qos = AsyncQueueSource_io_async_mem_5_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_id = AsyncQueueSource_io_async_mem_6_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_addr = AsyncQueueSource_io_async_mem_6_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_len = AsyncQueueSource_io_async_mem_6_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_size = AsyncQueueSource_io_async_mem_6_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_burst = AsyncQueueSource_io_async_mem_6_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_lock = AsyncQueueSource_io_async_mem_6_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_cache = AsyncQueueSource_io_async_mem_6_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_prot = AsyncQueueSource_io_async_mem_6_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_6_qos = AsyncQueueSource_io_async_mem_6_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_id = AsyncQueueSource_io_async_mem_7_id; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_addr = AsyncQueueSource_io_async_mem_7_addr; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_len = AsyncQueueSource_io_async_mem_7_len; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_size = AsyncQueueSource_io_async_mem_7_size; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_burst = AsyncQueueSource_io_async_mem_7_burst; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_lock = AsyncQueueSource_io_async_mem_7_lock; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_cache = AsyncQueueSource_io_async_mem_7_cache; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_prot = AsyncQueueSource_io_async_mem_7_prot; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_mem_7_qos = AsyncQueueSource_io_async_mem_7_qos; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_widx = AsyncQueueSource_io_async_widx; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_safe_widx_valid = AsyncQueueSource_io_async_safe_widx_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_ar_safe_source_reset_n = AsyncQueueSource_io_async_safe_source_reset_n; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_r_ridx = AsyncQueueSink_io_async_ridx; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_r_safe_ridx_valid = AsyncQueueSink_io_async_safe_ridx_valid; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign auto_out_r_safe_sink_reset_n = AsyncQueueSink_io_async_safe_sink_reset_n; // @[LazyModule.scala 173:49:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310699.4]
  assign AsyncQueueSource_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310702.4]
  assign AsyncQueueSource_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310703.4]
  assign AsyncQueueSource_io_enq_valid = auto_in_ar_valid; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310705.4]
  assign AsyncQueueSource_io_enq_bits_id = auto_in_ar_bits_id; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_enq_bits_addr = auto_in_ar_bits_addr; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_enq_bits_len = auto_in_ar_bits_len; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_enq_bits_size = auto_in_ar_bits_size; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_enq_bits_burst = auto_in_ar_bits_burst; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_enq_bits_lock = auto_in_ar_bits_lock; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_enq_bits_cache = auto_in_ar_bits_cache; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_enq_bits_prot = auto_in_ar_bits_prot; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_enq_bits_qos = auto_in_ar_bits_qos; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310704.4]
  assign AsyncQueueSource_io_async_ridx = auto_out_ar_ridx; // @[AsyncCrossing.scala 23:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310707.4]
  assign AsyncQueueSource_io_async_safe_ridx_valid = auto_out_ar_safe_ridx_valid; // @[AsyncCrossing.scala 23:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310707.4]
  assign AsyncQueueSource_io_async_safe_sink_reset_n = auto_out_ar_safe_sink_reset_n; // @[AsyncCrossing.scala 23:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310707.4]
  assign AsyncQueueSource_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310709.4]
  assign AsyncQueueSource_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310710.4]
  assign AsyncQueueSource_1_io_enq_valid = auto_in_aw_valid; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310712.4]
  assign AsyncQueueSource_1_io_enq_bits_id = auto_in_aw_bits_id; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_enq_bits_addr = auto_in_aw_bits_addr; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_enq_bits_len = auto_in_aw_bits_len; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_enq_bits_size = auto_in_aw_bits_size; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_enq_bits_burst = auto_in_aw_bits_burst; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_enq_bits_lock = auto_in_aw_bits_lock; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_enq_bits_cache = auto_in_aw_bits_cache; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_enq_bits_prot = auto_in_aw_bits_prot; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_enq_bits_qos = auto_in_aw_bits_qos; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310711.4]
  assign AsyncQueueSource_1_io_async_ridx = auto_out_aw_ridx; // @[AsyncCrossing.scala 24:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310714.4]
  assign AsyncQueueSource_1_io_async_safe_ridx_valid = auto_out_aw_safe_ridx_valid; // @[AsyncCrossing.scala 24:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310714.4]
  assign AsyncQueueSource_1_io_async_safe_sink_reset_n = auto_out_aw_safe_sink_reset_n; // @[AsyncCrossing.scala 24:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310714.4]
  assign AsyncQueueSource_2_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310716.4]
  assign AsyncQueueSource_2_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310717.4]
  assign AsyncQueueSource_2_io_enq_valid = auto_in_w_valid; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310719.4]
  assign AsyncQueueSource_2_io_enq_bits_data = auto_in_w_bits_data; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310718.4]
  assign AsyncQueueSource_2_io_enq_bits_strb = auto_in_w_bits_strb; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310718.4]
  assign AsyncQueueSource_2_io_enq_bits_last = auto_in_w_bits_last; // @[AsyncQueue.scala 193:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310718.4]
  assign AsyncQueueSource_2_io_async_ridx = auto_out_w_ridx; // @[AsyncCrossing.scala 25:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310721.4]
  assign AsyncQueueSource_2_io_async_safe_ridx_valid = auto_out_w_safe_ridx_valid; // @[AsyncCrossing.scala 25:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310721.4]
  assign AsyncQueueSource_2_io_async_safe_sink_reset_n = auto_out_w_safe_sink_reset_n; // @[AsyncCrossing.scala 25:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310721.4]
  assign AsyncQueueSink_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310723.4]
  assign AsyncQueueSink_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310724.4]
  assign AsyncQueueSink_io_deq_ready = auto_in_r_ready; // @[AsyncCrossing.scala 26:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310739.4]
  assign AsyncQueueSink_io_async_mem_0_id = auto_out_r_mem_0_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310731.4]
  assign AsyncQueueSink_io_async_mem_0_data = auto_out_r_mem_0_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310731.4]
  assign AsyncQueueSink_io_async_mem_0_resp = auto_out_r_mem_0_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310731.4]
  assign AsyncQueueSink_io_async_mem_0_last = auto_out_r_mem_0_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310731.4]
  assign AsyncQueueSink_io_async_mem_1_id = auto_out_r_mem_1_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310732.4]
  assign AsyncQueueSink_io_async_mem_1_data = auto_out_r_mem_1_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310732.4]
  assign AsyncQueueSink_io_async_mem_1_resp = auto_out_r_mem_1_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310732.4]
  assign AsyncQueueSink_io_async_mem_1_last = auto_out_r_mem_1_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310732.4]
  assign AsyncQueueSink_io_async_mem_2_id = auto_out_r_mem_2_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310733.4]
  assign AsyncQueueSink_io_async_mem_2_data = auto_out_r_mem_2_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310733.4]
  assign AsyncQueueSink_io_async_mem_2_resp = auto_out_r_mem_2_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310733.4]
  assign AsyncQueueSink_io_async_mem_2_last = auto_out_r_mem_2_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310733.4]
  assign AsyncQueueSink_io_async_mem_3_id = auto_out_r_mem_3_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310734.4]
  assign AsyncQueueSink_io_async_mem_3_data = auto_out_r_mem_3_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310734.4]
  assign AsyncQueueSink_io_async_mem_3_resp = auto_out_r_mem_3_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310734.4]
  assign AsyncQueueSink_io_async_mem_3_last = auto_out_r_mem_3_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310734.4]
  assign AsyncQueueSink_io_async_mem_4_id = auto_out_r_mem_4_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310735.4]
  assign AsyncQueueSink_io_async_mem_4_data = auto_out_r_mem_4_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310735.4]
  assign AsyncQueueSink_io_async_mem_4_resp = auto_out_r_mem_4_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310735.4]
  assign AsyncQueueSink_io_async_mem_4_last = auto_out_r_mem_4_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310735.4]
  assign AsyncQueueSink_io_async_mem_5_id = auto_out_r_mem_5_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310736.4]
  assign AsyncQueueSink_io_async_mem_5_data = auto_out_r_mem_5_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310736.4]
  assign AsyncQueueSink_io_async_mem_5_resp = auto_out_r_mem_5_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310736.4]
  assign AsyncQueueSink_io_async_mem_5_last = auto_out_r_mem_5_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310736.4]
  assign AsyncQueueSink_io_async_mem_6_id = auto_out_r_mem_6_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310737.4]
  assign AsyncQueueSink_io_async_mem_6_data = auto_out_r_mem_6_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310737.4]
  assign AsyncQueueSink_io_async_mem_6_resp = auto_out_r_mem_6_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310737.4]
  assign AsyncQueueSink_io_async_mem_6_last = auto_out_r_mem_6_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310737.4]
  assign AsyncQueueSink_io_async_mem_7_id = auto_out_r_mem_7_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310738.4]
  assign AsyncQueueSink_io_async_mem_7_data = auto_out_r_mem_7_data; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310738.4]
  assign AsyncQueueSink_io_async_mem_7_resp = auto_out_r_mem_7_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310738.4]
  assign AsyncQueueSink_io_async_mem_7_last = auto_out_r_mem_7_last; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310738.4]
  assign AsyncQueueSink_io_async_widx = auto_out_r_widx; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310729.4]
  assign AsyncQueueSink_io_async_safe_widx_valid = auto_out_r_safe_widx_valid; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310727.4]
  assign AsyncQueueSink_io_async_safe_source_reset_n = auto_out_r_safe_source_reset_n; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310726.4]
  assign AsyncQueueSink_1_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310741.4]
  assign AsyncQueueSink_1_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310742.4]
  assign AsyncQueueSink_1_io_deq_ready = auto_in_b_ready; // @[AsyncCrossing.scala 27:14:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310757.4]
  assign AsyncQueueSink_1_io_async_mem_0_id = auto_out_b_mem_0_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310749.4]
  assign AsyncQueueSink_1_io_async_mem_0_resp = auto_out_b_mem_0_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310749.4]
  assign AsyncQueueSink_1_io_async_mem_1_id = auto_out_b_mem_1_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310750.4]
  assign AsyncQueueSink_1_io_async_mem_1_resp = auto_out_b_mem_1_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310750.4]
  assign AsyncQueueSink_1_io_async_mem_2_id = auto_out_b_mem_2_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310751.4]
  assign AsyncQueueSink_1_io_async_mem_2_resp = auto_out_b_mem_2_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310751.4]
  assign AsyncQueueSink_1_io_async_mem_3_id = auto_out_b_mem_3_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310752.4]
  assign AsyncQueueSink_1_io_async_mem_3_resp = auto_out_b_mem_3_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310752.4]
  assign AsyncQueueSink_1_io_async_mem_4_id = auto_out_b_mem_4_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310753.4]
  assign AsyncQueueSink_1_io_async_mem_4_resp = auto_out_b_mem_4_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310753.4]
  assign AsyncQueueSink_1_io_async_mem_5_id = auto_out_b_mem_5_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310754.4]
  assign AsyncQueueSink_1_io_async_mem_5_resp = auto_out_b_mem_5_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310754.4]
  assign AsyncQueueSink_1_io_async_mem_6_id = auto_out_b_mem_6_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310755.4]
  assign AsyncQueueSink_1_io_async_mem_6_resp = auto_out_b_mem_6_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310755.4]
  assign AsyncQueueSink_1_io_async_mem_7_id = auto_out_b_mem_7_id; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310756.4]
  assign AsyncQueueSink_1_io_async_mem_7_resp = auto_out_b_mem_7_resp; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310756.4]
  assign AsyncQueueSink_1_io_async_widx = auto_out_b_widx; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310747.4]
  assign AsyncQueueSink_1_io_async_safe_widx_valid = auto_out_b_safe_widx_valid; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310745.4]
  assign AsyncQueueSink_1_io_async_safe_source_reset_n = auto_out_b_safe_source_reset_n; // @[AsyncQueue.scala 184:19:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310744.4]
endmodule
module XilinxVC707MIG( // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310759.2]
  input         clock, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310760.4]
  input         reset, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310761.4]
  output        auto_buffer_in_a_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  input         auto_buffer_in_a_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  input  [2:0]  auto_buffer_in_a_bits_opcode, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  input  [2:0]  auto_buffer_in_a_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  input  [6:0]  auto_buffer_in_a_bits_source, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  input  [31:0] auto_buffer_in_a_bits_address, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  input  [7:0]  auto_buffer_in_a_bits_mask, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  input  [63:0] auto_buffer_in_a_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  input         auto_buffer_in_d_ready, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output        auto_buffer_in_d_valid, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output [2:0]  auto_buffer_in_d_bits_opcode, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output [1:0]  auto_buffer_in_d_bits_param, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output [2:0]  auto_buffer_in_d_bits_size, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output [6:0]  auto_buffer_in_d_bits_source, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output        auto_buffer_in_d_bits_denied, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output [63:0] auto_buffer_in_d_bits_data, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output        auto_buffer_in_d_bits_corrupt, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310762.4]
  output [13:0] io_port_ddr3_addr, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output [2:0]  io_port_ddr3_ba, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_ras_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_cas_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_we_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_reset_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_ck_p, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_ck_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_cke, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_cs_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output [7:0]  io_port_ddr3_dm, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ddr3_odt, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  inout  [63:0] io_port_ddr3_dq, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  inout  [7:0]  io_port_ddr3_dqs_n, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  inout  [7:0]  io_port_ddr3_dqs_p, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  input         io_port_sys_clk_i, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ui_clk, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_ui_clk_sync_rst, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  output        io_port_mmcm_locked, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  input         io_port_aresetn, // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
  input         io_port_sys_rst // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310763.4]
);
  wire  buffer_clock; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_reset; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_in_a_ready; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_in_a_valid; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [2:0] buffer_auto_in_a_bits_size; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [6:0] buffer_auto_in_a_bits_source; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [31:0] buffer_auto_in_a_bits_address; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [63:0] buffer_auto_in_a_bits_data; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_in_d_ready; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_in_d_valid; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [1:0] buffer_auto_in_d_bits_param; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [2:0] buffer_auto_in_d_bits_size; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [6:0] buffer_auto_in_d_bits_source; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_in_d_bits_denied; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [63:0] buffer_auto_in_d_bits_data; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_in_d_bits_corrupt; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_out_a_ready; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_out_a_valid; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [2:0] buffer_auto_out_a_bits_size; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [6:0] buffer_auto_out_a_bits_source; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [31:0] buffer_auto_out_a_bits_address; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [63:0] buffer_auto_out_a_bits_data; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_out_d_ready; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_out_d_valid; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [2:0] buffer_auto_out_d_bits_size; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [6:0] buffer_auto_out_d_bits_source; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_out_d_bits_denied; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire [63:0] buffer_auto_out_d_bits_data; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  buffer_auto_out_d_bits_corrupt; // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
  wire  toaxi4_clock; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_reset; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_in_a_ready; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_in_a_valid; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [2:0] toaxi4_auto_in_a_bits_opcode; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [2:0] toaxi4_auto_in_a_bits_size; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [6:0] toaxi4_auto_in_a_bits_source; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [31:0] toaxi4_auto_in_a_bits_address; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [7:0] toaxi4_auto_in_a_bits_mask; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [63:0] toaxi4_auto_in_a_bits_data; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_in_d_ready; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_in_d_valid; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [2:0] toaxi4_auto_in_d_bits_opcode; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [2:0] toaxi4_auto_in_d_bits_size; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [6:0] toaxi4_auto_in_d_bits_source; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_in_d_bits_denied; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [63:0] toaxi4_auto_in_d_bits_data; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_in_d_bits_corrupt; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_aw_ready; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_aw_valid; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [5:0] toaxi4_auto_out_aw_bits_id; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [31:0] toaxi4_auto_out_aw_bits_addr; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [7:0] toaxi4_auto_out_aw_bits_len; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [2:0] toaxi4_auto_out_aw_bits_size; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [1:0] toaxi4_auto_out_aw_bits_burst; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_aw_bits_lock; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [3:0] toaxi4_auto_out_aw_bits_cache; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [2:0] toaxi4_auto_out_aw_bits_prot; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [3:0] toaxi4_auto_out_aw_bits_qos; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [10:0] toaxi4_auto_out_aw_bits_user; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_w_ready; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_w_valid; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [63:0] toaxi4_auto_out_w_bits_data; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [7:0] toaxi4_auto_out_w_bits_strb; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_w_bits_last; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_b_ready; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_b_valid; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [5:0] toaxi4_auto_out_b_bits_id; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [1:0] toaxi4_auto_out_b_bits_resp; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [10:0] toaxi4_auto_out_b_bits_user; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_ar_ready; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_ar_valid; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [5:0] toaxi4_auto_out_ar_bits_id; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [31:0] toaxi4_auto_out_ar_bits_addr; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [7:0] toaxi4_auto_out_ar_bits_len; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [2:0] toaxi4_auto_out_ar_bits_size; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [1:0] toaxi4_auto_out_ar_bits_burst; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_ar_bits_lock; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [3:0] toaxi4_auto_out_ar_bits_cache; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [2:0] toaxi4_auto_out_ar_bits_prot; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [3:0] toaxi4_auto_out_ar_bits_qos; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [10:0] toaxi4_auto_out_ar_bits_user; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_r_ready; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_r_valid; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [5:0] toaxi4_auto_out_r_bits_id; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [63:0] toaxi4_auto_out_r_bits_data; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [1:0] toaxi4_auto_out_r_bits_resp; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire [10:0] toaxi4_auto_out_r_bits_user; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  toaxi4_auto_out_r_bits_last; // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
  wire  indexer_auto_in_aw_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_aw_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [5:0] indexer_auto_in_aw_bits_id; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [31:0] indexer_auto_in_aw_bits_addr; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [7:0] indexer_auto_in_aw_bits_len; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [2:0] indexer_auto_in_aw_bits_size; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [1:0] indexer_auto_in_aw_bits_burst; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_aw_bits_lock; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_in_aw_bits_cache; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [2:0] indexer_auto_in_aw_bits_prot; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_in_aw_bits_qos; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [10:0] indexer_auto_in_aw_bits_user; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_w_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_w_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [63:0] indexer_auto_in_w_bits_data; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [7:0] indexer_auto_in_w_bits_strb; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_w_bits_last; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_b_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_b_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [5:0] indexer_auto_in_b_bits_id; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [1:0] indexer_auto_in_b_bits_resp; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [10:0] indexer_auto_in_b_bits_user; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_ar_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_ar_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [5:0] indexer_auto_in_ar_bits_id; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [31:0] indexer_auto_in_ar_bits_addr; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [7:0] indexer_auto_in_ar_bits_len; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [2:0] indexer_auto_in_ar_bits_size; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [1:0] indexer_auto_in_ar_bits_burst; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_ar_bits_lock; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_in_ar_bits_cache; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [2:0] indexer_auto_in_ar_bits_prot; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_in_ar_bits_qos; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [10:0] indexer_auto_in_ar_bits_user; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_r_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_r_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [5:0] indexer_auto_in_r_bits_id; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [63:0] indexer_auto_in_r_bits_data; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [1:0] indexer_auto_in_r_bits_resp; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [10:0] indexer_auto_in_r_bits_user; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_in_r_bits_last; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_aw_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_aw_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_out_aw_bits_id; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [31:0] indexer_auto_out_aw_bits_addr; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [7:0] indexer_auto_out_aw_bits_len; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [2:0] indexer_auto_out_aw_bits_size; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [1:0] indexer_auto_out_aw_bits_burst; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_aw_bits_lock; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_out_aw_bits_cache; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [2:0] indexer_auto_out_aw_bits_prot; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_out_aw_bits_qos; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [12:0] indexer_auto_out_aw_bits_user; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_w_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_w_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [63:0] indexer_auto_out_w_bits_data; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [7:0] indexer_auto_out_w_bits_strb; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_w_bits_last; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_b_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_b_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_out_b_bits_id; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [1:0] indexer_auto_out_b_bits_resp; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [12:0] indexer_auto_out_b_bits_user; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_ar_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_ar_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_out_ar_bits_id; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [31:0] indexer_auto_out_ar_bits_addr; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [7:0] indexer_auto_out_ar_bits_len; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [2:0] indexer_auto_out_ar_bits_size; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [1:0] indexer_auto_out_ar_bits_burst; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_ar_bits_lock; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_out_ar_bits_cache; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [2:0] indexer_auto_out_ar_bits_prot; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_out_ar_bits_qos; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [12:0] indexer_auto_out_ar_bits_user; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_r_ready; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_r_valid; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [3:0] indexer_auto_out_r_bits_id; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [63:0] indexer_auto_out_r_bits_data; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [1:0] indexer_auto_out_r_bits_resp; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire [12:0] indexer_auto_out_r_bits_user; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  indexer_auto_out_r_bits_last; // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
  wire  deint_clock; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_reset; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_aw_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_aw_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_in_aw_bits_id; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [31:0] deint_auto_in_aw_bits_addr; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [7:0] deint_auto_in_aw_bits_len; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [2:0] deint_auto_in_aw_bits_size; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [1:0] deint_auto_in_aw_bits_burst; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_aw_bits_lock; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_in_aw_bits_cache; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [2:0] deint_auto_in_aw_bits_prot; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_in_aw_bits_qos; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [12:0] deint_auto_in_aw_bits_user; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_w_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_w_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [63:0] deint_auto_in_w_bits_data; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [7:0] deint_auto_in_w_bits_strb; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_w_bits_last; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_b_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_b_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_in_b_bits_id; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [1:0] deint_auto_in_b_bits_resp; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [12:0] deint_auto_in_b_bits_user; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_ar_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_ar_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_in_ar_bits_id; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [31:0] deint_auto_in_ar_bits_addr; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [7:0] deint_auto_in_ar_bits_len; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [2:0] deint_auto_in_ar_bits_size; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [1:0] deint_auto_in_ar_bits_burst; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_ar_bits_lock; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_in_ar_bits_cache; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [2:0] deint_auto_in_ar_bits_prot; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_in_ar_bits_qos; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [12:0] deint_auto_in_ar_bits_user; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_r_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_r_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_in_r_bits_id; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [63:0] deint_auto_in_r_bits_data; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [1:0] deint_auto_in_r_bits_resp; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [12:0] deint_auto_in_r_bits_user; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_in_r_bits_last; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_aw_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_aw_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_out_aw_bits_id; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [31:0] deint_auto_out_aw_bits_addr; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [7:0] deint_auto_out_aw_bits_len; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [2:0] deint_auto_out_aw_bits_size; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [1:0] deint_auto_out_aw_bits_burst; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_aw_bits_lock; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_out_aw_bits_cache; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [2:0] deint_auto_out_aw_bits_prot; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_out_aw_bits_qos; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [12:0] deint_auto_out_aw_bits_user; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_w_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_w_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [63:0] deint_auto_out_w_bits_data; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [7:0] deint_auto_out_w_bits_strb; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_w_bits_last; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_b_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_b_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_out_b_bits_id; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [1:0] deint_auto_out_b_bits_resp; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [12:0] deint_auto_out_b_bits_user; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_ar_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_ar_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_out_ar_bits_id; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [31:0] deint_auto_out_ar_bits_addr; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [7:0] deint_auto_out_ar_bits_len; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [2:0] deint_auto_out_ar_bits_size; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [1:0] deint_auto_out_ar_bits_burst; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_ar_bits_lock; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_out_ar_bits_cache; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [2:0] deint_auto_out_ar_bits_prot; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_out_ar_bits_qos; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [12:0] deint_auto_out_ar_bits_user; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_r_ready; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_r_valid; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [3:0] deint_auto_out_r_bits_id; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [63:0] deint_auto_out_r_bits_data; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [1:0] deint_auto_out_r_bits_resp; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire [12:0] deint_auto_out_r_bits_user; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  deint_auto_out_r_bits_last; // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
  wire  yank_clock; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_reset; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_aw_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_aw_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_in_aw_bits_id; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [31:0] yank_auto_in_aw_bits_addr; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [7:0] yank_auto_in_aw_bits_len; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [2:0] yank_auto_in_aw_bits_size; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [1:0] yank_auto_in_aw_bits_burst; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_aw_bits_lock; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_in_aw_bits_cache; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [2:0] yank_auto_in_aw_bits_prot; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_in_aw_bits_qos; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [12:0] yank_auto_in_aw_bits_user; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_w_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_w_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [63:0] yank_auto_in_w_bits_data; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [7:0] yank_auto_in_w_bits_strb; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_w_bits_last; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_b_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_b_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_in_b_bits_id; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [1:0] yank_auto_in_b_bits_resp; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [12:0] yank_auto_in_b_bits_user; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_ar_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_ar_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_in_ar_bits_id; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [31:0] yank_auto_in_ar_bits_addr; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [7:0] yank_auto_in_ar_bits_len; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [2:0] yank_auto_in_ar_bits_size; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [1:0] yank_auto_in_ar_bits_burst; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_ar_bits_lock; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_in_ar_bits_cache; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [2:0] yank_auto_in_ar_bits_prot; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_in_ar_bits_qos; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [12:0] yank_auto_in_ar_bits_user; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_r_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_r_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_in_r_bits_id; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [63:0] yank_auto_in_r_bits_data; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [1:0] yank_auto_in_r_bits_resp; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [12:0] yank_auto_in_r_bits_user; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_in_r_bits_last; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_aw_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_aw_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_out_aw_bits_id; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [31:0] yank_auto_out_aw_bits_addr; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [7:0] yank_auto_out_aw_bits_len; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [2:0] yank_auto_out_aw_bits_size; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [1:0] yank_auto_out_aw_bits_burst; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_aw_bits_lock; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_out_aw_bits_cache; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [2:0] yank_auto_out_aw_bits_prot; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_out_aw_bits_qos; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_w_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_w_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [63:0] yank_auto_out_w_bits_data; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [7:0] yank_auto_out_w_bits_strb; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_w_bits_last; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_b_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_b_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_out_b_bits_id; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [1:0] yank_auto_out_b_bits_resp; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_ar_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_ar_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_out_ar_bits_id; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [31:0] yank_auto_out_ar_bits_addr; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [7:0] yank_auto_out_ar_bits_len; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [2:0] yank_auto_out_ar_bits_size; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [1:0] yank_auto_out_ar_bits_burst; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_ar_bits_lock; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_out_ar_bits_cache; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [2:0] yank_auto_out_ar_bits_prot; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_out_ar_bits_qos; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_r_ready; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_r_valid; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] yank_auto_out_r_bits_id; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [63:0] yank_auto_out_r_bits_data; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [1:0] yank_auto_out_r_bits_resp; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire  yank_auto_out_r_bits_last; // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_0_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_aw_mem_0_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_aw_mem_0_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_0_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_aw_mem_0_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_mem_0_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_0_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_0_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_0_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_1_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_aw_mem_1_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_aw_mem_1_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_1_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_aw_mem_1_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_mem_1_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_1_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_1_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_1_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_2_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_aw_mem_2_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_aw_mem_2_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_2_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_aw_mem_2_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_mem_2_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_2_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_2_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_2_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_3_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_aw_mem_3_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_aw_mem_3_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_3_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_aw_mem_3_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_mem_3_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_3_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_3_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_3_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_4_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_aw_mem_4_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_aw_mem_4_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_4_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_aw_mem_4_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_mem_4_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_4_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_4_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_4_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_5_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_aw_mem_5_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_aw_mem_5_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_5_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_aw_mem_5_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_mem_5_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_5_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_5_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_5_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_6_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_aw_mem_6_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_aw_mem_6_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_6_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_aw_mem_6_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_mem_6_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_6_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_6_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_6_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_7_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_aw_mem_7_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_aw_mem_7_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_7_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_aw_mem_7_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_mem_7_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_7_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_aw_mem_7_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_mem_7_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_ridx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_aw_widx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_safe_ridx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_safe_widx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_safe_source_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_aw_safe_sink_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_w_mem_0_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_w_mem_0_strb; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_mem_0_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_w_mem_1_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_w_mem_1_strb; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_mem_1_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_w_mem_2_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_w_mem_2_strb; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_mem_2_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_w_mem_3_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_w_mem_3_strb; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_mem_3_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_w_mem_4_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_w_mem_4_strb; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_mem_4_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_w_mem_5_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_w_mem_5_strb; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_mem_5_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_w_mem_6_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_w_mem_6_strb; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_mem_6_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_w_mem_7_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_w_mem_7_strb; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_mem_7_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_w_ridx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_w_widx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_safe_ridx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_safe_widx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_safe_source_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_w_safe_sink_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_mem_0_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_b_mem_0_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_mem_1_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_b_mem_1_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_mem_2_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_b_mem_2_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_mem_3_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_b_mem_3_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_mem_4_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_b_mem_4_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_mem_5_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_b_mem_5_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_mem_6_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_b_mem_6_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_mem_7_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_b_mem_7_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_ridx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_b_widx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_b_safe_ridx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_b_safe_widx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_b_safe_source_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_b_safe_sink_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_0_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_ar_mem_0_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_ar_mem_0_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_0_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_ar_mem_0_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_mem_0_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_0_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_0_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_0_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_1_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_ar_mem_1_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_ar_mem_1_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_1_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_ar_mem_1_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_mem_1_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_1_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_1_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_1_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_2_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_ar_mem_2_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_ar_mem_2_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_2_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_ar_mem_2_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_mem_2_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_2_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_2_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_2_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_3_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_ar_mem_3_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_ar_mem_3_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_3_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_ar_mem_3_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_mem_3_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_3_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_3_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_3_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_4_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_ar_mem_4_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_ar_mem_4_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_4_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_ar_mem_4_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_mem_4_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_4_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_4_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_4_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_5_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_ar_mem_5_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_ar_mem_5_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_5_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_ar_mem_5_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_mem_5_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_5_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_5_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_5_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_6_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_ar_mem_6_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_ar_mem_6_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_6_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_ar_mem_6_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_mem_6_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_6_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_6_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_6_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_7_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [31:0] island_auto_axi4in_xing_in_ar_mem_7_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_auto_axi4in_xing_in_ar_mem_7_len; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_7_size; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_ar_mem_7_burst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_mem_7_lock; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_7_cache; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_auto_axi4in_xing_in_ar_mem_7_prot; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_mem_7_qos; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_ridx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_ar_widx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_safe_ridx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_safe_widx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_safe_source_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_ar_safe_sink_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_mem_0_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_r_mem_0_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_r_mem_0_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_mem_0_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_mem_1_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_r_mem_1_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_r_mem_1_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_mem_1_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_mem_2_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_r_mem_2_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_r_mem_2_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_mem_2_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_mem_3_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_r_mem_3_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_r_mem_3_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_mem_3_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_mem_4_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_r_mem_4_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_r_mem_4_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_mem_4_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_mem_5_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_r_mem_5_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_r_mem_5_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_mem_5_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_mem_6_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_r_mem_6_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_r_mem_6_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_mem_6_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_mem_7_id; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [63:0] island_auto_axi4in_xing_in_r_mem_7_data; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [1:0] island_auto_axi4in_xing_in_r_mem_7_resp; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_mem_7_last; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_ridx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [3:0] island_auto_axi4in_xing_in_r_widx; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_safe_ridx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_safe_widx_valid; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_safe_source_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_auto_axi4in_xing_in_r_safe_sink_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [13:0] island_io_port_ddr3_addr; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [2:0] island_io_port_ddr3_ba; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_ras_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_cas_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_we_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_reset_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_ck_p; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_ck_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_cke; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_cs_n; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire [7:0] island_io_port_ddr3_dm; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ddr3_odt; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_sys_clk_i; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ui_clk; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_ui_clk_sync_rst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_mmcm_locked; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_aresetn; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  island_io_port_sys_rst; // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
  wire  axi4asource_clock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_reset; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_aw_ready; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_aw_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_in_aw_bits_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_in_aw_bits_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_in_aw_bits_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_in_aw_bits_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_in_aw_bits_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_aw_bits_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_in_aw_bits_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_in_aw_bits_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_in_aw_bits_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_w_ready; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_w_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_in_w_bits_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_in_w_bits_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_w_bits_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_b_ready; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_b_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_in_b_bits_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_in_b_bits_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_ar_ready; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_ar_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_in_ar_bits_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_in_ar_bits_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_in_ar_bits_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_in_ar_bits_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_in_ar_bits_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_ar_bits_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_in_ar_bits_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_in_ar_bits_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_in_ar_bits_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_r_ready; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_r_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_in_r_bits_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_in_r_bits_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_in_r_bits_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_in_r_bits_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_0_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_aw_mem_0_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_aw_mem_0_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_0_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_aw_mem_0_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_mem_0_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_0_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_0_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_0_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_1_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_aw_mem_1_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_aw_mem_1_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_1_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_aw_mem_1_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_mem_1_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_1_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_1_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_1_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_2_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_aw_mem_2_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_aw_mem_2_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_2_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_aw_mem_2_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_mem_2_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_2_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_2_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_2_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_3_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_aw_mem_3_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_aw_mem_3_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_3_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_aw_mem_3_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_mem_3_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_3_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_3_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_3_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_4_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_aw_mem_4_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_aw_mem_4_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_4_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_aw_mem_4_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_mem_4_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_4_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_4_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_4_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_5_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_aw_mem_5_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_aw_mem_5_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_5_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_aw_mem_5_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_mem_5_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_5_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_5_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_5_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_6_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_aw_mem_6_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_aw_mem_6_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_6_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_aw_mem_6_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_mem_6_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_6_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_6_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_6_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_7_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_aw_mem_7_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_aw_mem_7_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_7_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_aw_mem_7_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_mem_7_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_7_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_aw_mem_7_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_mem_7_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_ridx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_aw_widx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_safe_ridx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_safe_widx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_safe_source_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_aw_safe_sink_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_w_mem_0_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_w_mem_0_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_mem_0_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_w_mem_1_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_w_mem_1_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_mem_1_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_w_mem_2_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_w_mem_2_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_mem_2_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_w_mem_3_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_w_mem_3_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_mem_3_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_w_mem_4_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_w_mem_4_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_mem_4_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_w_mem_5_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_w_mem_5_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_mem_5_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_w_mem_6_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_w_mem_6_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_mem_6_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_w_mem_7_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_w_mem_7_strb; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_mem_7_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_w_ridx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_w_widx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_safe_ridx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_safe_widx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_safe_source_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_w_safe_sink_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_mem_0_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_b_mem_0_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_mem_1_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_b_mem_1_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_mem_2_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_b_mem_2_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_mem_3_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_b_mem_3_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_mem_4_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_b_mem_4_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_mem_5_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_b_mem_5_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_mem_6_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_b_mem_6_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_mem_7_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_b_mem_7_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_ridx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_b_widx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_b_safe_ridx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_b_safe_widx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_b_safe_source_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_b_safe_sink_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_0_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_ar_mem_0_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_ar_mem_0_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_0_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_ar_mem_0_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_mem_0_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_0_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_0_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_0_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_1_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_ar_mem_1_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_ar_mem_1_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_1_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_ar_mem_1_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_mem_1_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_1_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_1_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_1_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_2_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_ar_mem_2_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_ar_mem_2_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_2_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_ar_mem_2_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_mem_2_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_2_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_2_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_2_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_3_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_ar_mem_3_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_ar_mem_3_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_3_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_ar_mem_3_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_mem_3_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_3_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_3_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_3_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_4_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_ar_mem_4_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_ar_mem_4_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_4_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_ar_mem_4_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_mem_4_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_4_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_4_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_4_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_5_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_ar_mem_5_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_ar_mem_5_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_5_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_ar_mem_5_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_mem_5_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_5_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_5_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_5_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_6_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_ar_mem_6_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_ar_mem_6_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_6_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_ar_mem_6_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_mem_6_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_6_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_6_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_6_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_7_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [31:0] axi4asource_auto_out_ar_mem_7_addr; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [7:0] axi4asource_auto_out_ar_mem_7_len; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_7_size; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_ar_mem_7_burst; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_mem_7_lock; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_7_cache; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [2:0] axi4asource_auto_out_ar_mem_7_prot; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_mem_7_qos; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_ridx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_ar_widx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_safe_ridx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_safe_widx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_safe_source_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_ar_safe_sink_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_mem_0_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_r_mem_0_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_r_mem_0_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_mem_0_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_mem_1_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_r_mem_1_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_r_mem_1_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_mem_1_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_mem_2_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_r_mem_2_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_r_mem_2_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_mem_2_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_mem_3_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_r_mem_3_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_r_mem_3_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_mem_3_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_mem_4_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_r_mem_4_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_r_mem_4_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_mem_4_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_mem_5_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_r_mem_5_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_r_mem_5_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_mem_5_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_mem_6_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_r_mem_6_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_r_mem_6_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_mem_6_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_mem_7_id; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [63:0] axi4asource_auto_out_r_mem_7_data; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [1:0] axi4asource_auto_out_r_mem_7_resp; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_mem_7_last; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_ridx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire [3:0] axi4asource_auto_out_r_widx; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_safe_ridx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_safe_widx_valid; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_safe_source_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  wire  axi4asource_auto_out_r_safe_sink_reset_n; // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
  TLBuffer_33 buffer ( // @[XilinxVC707MIG.scala 153:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310769.4]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
  );
  TLToAXI4 toaxi4 ( // @[XilinxVC707MIG.scala 154:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310775.4]
    .clock(toaxi4_clock),
    .reset(toaxi4_reset),
    .auto_in_a_ready(toaxi4_auto_in_a_ready),
    .auto_in_a_valid(toaxi4_auto_in_a_valid),
    .auto_in_a_bits_opcode(toaxi4_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(toaxi4_auto_in_a_bits_size),
    .auto_in_a_bits_source(toaxi4_auto_in_a_bits_source),
    .auto_in_a_bits_address(toaxi4_auto_in_a_bits_address),
    .auto_in_a_bits_mask(toaxi4_auto_in_a_bits_mask),
    .auto_in_a_bits_data(toaxi4_auto_in_a_bits_data),
    .auto_in_d_ready(toaxi4_auto_in_d_ready),
    .auto_in_d_valid(toaxi4_auto_in_d_valid),
    .auto_in_d_bits_opcode(toaxi4_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(toaxi4_auto_in_d_bits_size),
    .auto_in_d_bits_source(toaxi4_auto_in_d_bits_source),
    .auto_in_d_bits_denied(toaxi4_auto_in_d_bits_denied),
    .auto_in_d_bits_data(toaxi4_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(toaxi4_auto_in_d_bits_corrupt),
    .auto_out_aw_ready(toaxi4_auto_out_aw_ready),
    .auto_out_aw_valid(toaxi4_auto_out_aw_valid),
    .auto_out_aw_bits_id(toaxi4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(toaxi4_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(toaxi4_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(toaxi4_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(toaxi4_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(toaxi4_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(toaxi4_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(toaxi4_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(toaxi4_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(toaxi4_auto_out_aw_bits_user),
    .auto_out_w_ready(toaxi4_auto_out_w_ready),
    .auto_out_w_valid(toaxi4_auto_out_w_valid),
    .auto_out_w_bits_data(toaxi4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(toaxi4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(toaxi4_auto_out_w_bits_last),
    .auto_out_b_ready(toaxi4_auto_out_b_ready),
    .auto_out_b_valid(toaxi4_auto_out_b_valid),
    .auto_out_b_bits_id(toaxi4_auto_out_b_bits_id),
    .auto_out_b_bits_resp(toaxi4_auto_out_b_bits_resp),
    .auto_out_b_bits_user(toaxi4_auto_out_b_bits_user),
    .auto_out_ar_ready(toaxi4_auto_out_ar_ready),
    .auto_out_ar_valid(toaxi4_auto_out_ar_valid),
    .auto_out_ar_bits_id(toaxi4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(toaxi4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(toaxi4_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(toaxi4_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(toaxi4_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(toaxi4_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(toaxi4_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(toaxi4_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(toaxi4_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(toaxi4_auto_out_ar_bits_user),
    .auto_out_r_ready(toaxi4_auto_out_r_ready),
    .auto_out_r_valid(toaxi4_auto_out_r_valid),
    .auto_out_r_bits_id(toaxi4_auto_out_r_bits_id),
    .auto_out_r_bits_data(toaxi4_auto_out_r_bits_data),
    .auto_out_r_bits_resp(toaxi4_auto_out_r_bits_resp),
    .auto_out_r_bits_user(toaxi4_auto_out_r_bits_user),
    .auto_out_r_bits_last(toaxi4_auto_out_r_bits_last)
  );
  AXI4IdIndexer indexer ( // @[XilinxVC707MIG.scala 155:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310781.4]
    .auto_in_aw_ready(indexer_auto_in_aw_ready),
    .auto_in_aw_valid(indexer_auto_in_aw_valid),
    .auto_in_aw_bits_id(indexer_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(indexer_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(indexer_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(indexer_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(indexer_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(indexer_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(indexer_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(indexer_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(indexer_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(indexer_auto_in_aw_bits_user),
    .auto_in_w_ready(indexer_auto_in_w_ready),
    .auto_in_w_valid(indexer_auto_in_w_valid),
    .auto_in_w_bits_data(indexer_auto_in_w_bits_data),
    .auto_in_w_bits_strb(indexer_auto_in_w_bits_strb),
    .auto_in_w_bits_last(indexer_auto_in_w_bits_last),
    .auto_in_b_ready(indexer_auto_in_b_ready),
    .auto_in_b_valid(indexer_auto_in_b_valid),
    .auto_in_b_bits_id(indexer_auto_in_b_bits_id),
    .auto_in_b_bits_resp(indexer_auto_in_b_bits_resp),
    .auto_in_b_bits_user(indexer_auto_in_b_bits_user),
    .auto_in_ar_ready(indexer_auto_in_ar_ready),
    .auto_in_ar_valid(indexer_auto_in_ar_valid),
    .auto_in_ar_bits_id(indexer_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(indexer_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(indexer_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(indexer_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(indexer_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(indexer_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(indexer_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(indexer_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(indexer_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(indexer_auto_in_ar_bits_user),
    .auto_in_r_ready(indexer_auto_in_r_ready),
    .auto_in_r_valid(indexer_auto_in_r_valid),
    .auto_in_r_bits_id(indexer_auto_in_r_bits_id),
    .auto_in_r_bits_data(indexer_auto_in_r_bits_data),
    .auto_in_r_bits_resp(indexer_auto_in_r_bits_resp),
    .auto_in_r_bits_user(indexer_auto_in_r_bits_user),
    .auto_in_r_bits_last(indexer_auto_in_r_bits_last),
    .auto_out_aw_ready(indexer_auto_out_aw_ready),
    .auto_out_aw_valid(indexer_auto_out_aw_valid),
    .auto_out_aw_bits_id(indexer_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(indexer_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(indexer_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(indexer_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(indexer_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(indexer_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(indexer_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(indexer_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(indexer_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(indexer_auto_out_aw_bits_user),
    .auto_out_w_ready(indexer_auto_out_w_ready),
    .auto_out_w_valid(indexer_auto_out_w_valid),
    .auto_out_w_bits_data(indexer_auto_out_w_bits_data),
    .auto_out_w_bits_strb(indexer_auto_out_w_bits_strb),
    .auto_out_w_bits_last(indexer_auto_out_w_bits_last),
    .auto_out_b_ready(indexer_auto_out_b_ready),
    .auto_out_b_valid(indexer_auto_out_b_valid),
    .auto_out_b_bits_id(indexer_auto_out_b_bits_id),
    .auto_out_b_bits_resp(indexer_auto_out_b_bits_resp),
    .auto_out_b_bits_user(indexer_auto_out_b_bits_user),
    .auto_out_ar_ready(indexer_auto_out_ar_ready),
    .auto_out_ar_valid(indexer_auto_out_ar_valid),
    .auto_out_ar_bits_id(indexer_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(indexer_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(indexer_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(indexer_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(indexer_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(indexer_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(indexer_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(indexer_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(indexer_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(indexer_auto_out_ar_bits_user),
    .auto_out_r_ready(indexer_auto_out_r_ready),
    .auto_out_r_valid(indexer_auto_out_r_valid),
    .auto_out_r_bits_id(indexer_auto_out_r_bits_id),
    .auto_out_r_bits_data(indexer_auto_out_r_bits_data),
    .auto_out_r_bits_resp(indexer_auto_out_r_bits_resp),
    .auto_out_r_bits_user(indexer_auto_out_r_bits_user),
    .auto_out_r_bits_last(indexer_auto_out_r_bits_last)
  );
  AXI4Deinterleaver deint ( // @[XilinxVC707MIG.scala 156:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310787.4]
    .clock(deint_clock),
    .reset(deint_reset),
    .auto_in_aw_ready(deint_auto_in_aw_ready),
    .auto_in_aw_valid(deint_auto_in_aw_valid),
    .auto_in_aw_bits_id(deint_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(deint_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(deint_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(deint_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(deint_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(deint_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(deint_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(deint_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(deint_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(deint_auto_in_aw_bits_user),
    .auto_in_w_ready(deint_auto_in_w_ready),
    .auto_in_w_valid(deint_auto_in_w_valid),
    .auto_in_w_bits_data(deint_auto_in_w_bits_data),
    .auto_in_w_bits_strb(deint_auto_in_w_bits_strb),
    .auto_in_w_bits_last(deint_auto_in_w_bits_last),
    .auto_in_b_ready(deint_auto_in_b_ready),
    .auto_in_b_valid(deint_auto_in_b_valid),
    .auto_in_b_bits_id(deint_auto_in_b_bits_id),
    .auto_in_b_bits_resp(deint_auto_in_b_bits_resp),
    .auto_in_b_bits_user(deint_auto_in_b_bits_user),
    .auto_in_ar_ready(deint_auto_in_ar_ready),
    .auto_in_ar_valid(deint_auto_in_ar_valid),
    .auto_in_ar_bits_id(deint_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(deint_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(deint_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(deint_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(deint_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(deint_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(deint_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(deint_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(deint_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(deint_auto_in_ar_bits_user),
    .auto_in_r_ready(deint_auto_in_r_ready),
    .auto_in_r_valid(deint_auto_in_r_valid),
    .auto_in_r_bits_id(deint_auto_in_r_bits_id),
    .auto_in_r_bits_data(deint_auto_in_r_bits_data),
    .auto_in_r_bits_resp(deint_auto_in_r_bits_resp),
    .auto_in_r_bits_user(deint_auto_in_r_bits_user),
    .auto_in_r_bits_last(deint_auto_in_r_bits_last),
    .auto_out_aw_ready(deint_auto_out_aw_ready),
    .auto_out_aw_valid(deint_auto_out_aw_valid),
    .auto_out_aw_bits_id(deint_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(deint_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(deint_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(deint_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(deint_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(deint_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(deint_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(deint_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(deint_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(deint_auto_out_aw_bits_user),
    .auto_out_w_ready(deint_auto_out_w_ready),
    .auto_out_w_valid(deint_auto_out_w_valid),
    .auto_out_w_bits_data(deint_auto_out_w_bits_data),
    .auto_out_w_bits_strb(deint_auto_out_w_bits_strb),
    .auto_out_w_bits_last(deint_auto_out_w_bits_last),
    .auto_out_b_ready(deint_auto_out_b_ready),
    .auto_out_b_valid(deint_auto_out_b_valid),
    .auto_out_b_bits_id(deint_auto_out_b_bits_id),
    .auto_out_b_bits_resp(deint_auto_out_b_bits_resp),
    .auto_out_b_bits_user(deint_auto_out_b_bits_user),
    .auto_out_ar_ready(deint_auto_out_ar_ready),
    .auto_out_ar_valid(deint_auto_out_ar_valid),
    .auto_out_ar_bits_id(deint_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(deint_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(deint_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(deint_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(deint_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(deint_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(deint_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(deint_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(deint_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(deint_auto_out_ar_bits_user),
    .auto_out_r_ready(deint_auto_out_r_ready),
    .auto_out_r_valid(deint_auto_out_r_valid),
    .auto_out_r_bits_id(deint_auto_out_r_bits_id),
    .auto_out_r_bits_data(deint_auto_out_r_bits_data),
    .auto_out_r_bits_resp(deint_auto_out_r_bits_resp),
    .auto_out_r_bits_user(deint_auto_out_r_bits_user),
    .auto_out_r_bits_last(deint_auto_out_r_bits_last)
  );
  AXI4UserYanker yank ( // @[XilinxVC707MIG.scala 157:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310793.4]
    .clock(yank_clock),
    .reset(yank_reset),
    .auto_in_aw_ready(yank_auto_in_aw_ready),
    .auto_in_aw_valid(yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(yank_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(yank_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(yank_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(yank_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(yank_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(yank_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(yank_auto_in_aw_bits_user),
    .auto_in_w_ready(yank_auto_in_w_ready),
    .auto_in_w_valid(yank_auto_in_w_valid),
    .auto_in_w_bits_data(yank_auto_in_w_bits_data),
    .auto_in_w_bits_strb(yank_auto_in_w_bits_strb),
    .auto_in_w_bits_last(yank_auto_in_w_bits_last),
    .auto_in_b_ready(yank_auto_in_b_ready),
    .auto_in_b_valid(yank_auto_in_b_valid),
    .auto_in_b_bits_id(yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(yank_auto_in_b_bits_resp),
    .auto_in_b_bits_user(yank_auto_in_b_bits_user),
    .auto_in_ar_ready(yank_auto_in_ar_ready),
    .auto_in_ar_valid(yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(yank_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(yank_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(yank_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(yank_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(yank_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(yank_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(yank_auto_in_ar_bits_user),
    .auto_in_r_ready(yank_auto_in_r_ready),
    .auto_in_r_valid(yank_auto_in_r_valid),
    .auto_in_r_bits_id(yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(yank_auto_in_r_bits_resp),
    .auto_in_r_bits_user(yank_auto_in_r_bits_user),
    .auto_in_r_bits_last(yank_auto_in_r_bits_last),
    .auto_out_aw_ready(yank_auto_out_aw_ready),
    .auto_out_aw_valid(yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(yank_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(yank_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(yank_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(yank_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(yank_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(yank_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(yank_auto_out_aw_bits_qos),
    .auto_out_w_ready(yank_auto_out_w_ready),
    .auto_out_w_valid(yank_auto_out_w_valid),
    .auto_out_w_bits_data(yank_auto_out_w_bits_data),
    .auto_out_w_bits_strb(yank_auto_out_w_bits_strb),
    .auto_out_w_bits_last(yank_auto_out_w_bits_last),
    .auto_out_b_ready(yank_auto_out_b_ready),
    .auto_out_b_valid(yank_auto_out_b_valid),
    .auto_out_b_bits_id(yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(yank_auto_out_ar_ready),
    .auto_out_ar_valid(yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(yank_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(yank_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(yank_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(yank_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(yank_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(yank_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(yank_auto_out_ar_bits_qos),
    .auto_out_r_ready(yank_auto_out_r_ready),
    .auto_out_r_valid(yank_auto_out_r_valid),
    .auto_out_r_bits_id(yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(yank_auto_out_r_bits_last)
  );
  XilinxVC707MIGIsland island ( // @[XilinxVC707MIG.scala 158:27:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310799.4]
    .auto_axi4in_xing_in_aw_mem_0_id(island_auto_axi4in_xing_in_aw_mem_0_id),
    .auto_axi4in_xing_in_aw_mem_0_addr(island_auto_axi4in_xing_in_aw_mem_0_addr),
    .auto_axi4in_xing_in_aw_mem_0_len(island_auto_axi4in_xing_in_aw_mem_0_len),
    .auto_axi4in_xing_in_aw_mem_0_size(island_auto_axi4in_xing_in_aw_mem_0_size),
    .auto_axi4in_xing_in_aw_mem_0_burst(island_auto_axi4in_xing_in_aw_mem_0_burst),
    .auto_axi4in_xing_in_aw_mem_0_lock(island_auto_axi4in_xing_in_aw_mem_0_lock),
    .auto_axi4in_xing_in_aw_mem_0_cache(island_auto_axi4in_xing_in_aw_mem_0_cache),
    .auto_axi4in_xing_in_aw_mem_0_prot(island_auto_axi4in_xing_in_aw_mem_0_prot),
    .auto_axi4in_xing_in_aw_mem_0_qos(island_auto_axi4in_xing_in_aw_mem_0_qos),
    .auto_axi4in_xing_in_aw_mem_1_id(island_auto_axi4in_xing_in_aw_mem_1_id),
    .auto_axi4in_xing_in_aw_mem_1_addr(island_auto_axi4in_xing_in_aw_mem_1_addr),
    .auto_axi4in_xing_in_aw_mem_1_len(island_auto_axi4in_xing_in_aw_mem_1_len),
    .auto_axi4in_xing_in_aw_mem_1_size(island_auto_axi4in_xing_in_aw_mem_1_size),
    .auto_axi4in_xing_in_aw_mem_1_burst(island_auto_axi4in_xing_in_aw_mem_1_burst),
    .auto_axi4in_xing_in_aw_mem_1_lock(island_auto_axi4in_xing_in_aw_mem_1_lock),
    .auto_axi4in_xing_in_aw_mem_1_cache(island_auto_axi4in_xing_in_aw_mem_1_cache),
    .auto_axi4in_xing_in_aw_mem_1_prot(island_auto_axi4in_xing_in_aw_mem_1_prot),
    .auto_axi4in_xing_in_aw_mem_1_qos(island_auto_axi4in_xing_in_aw_mem_1_qos),
    .auto_axi4in_xing_in_aw_mem_2_id(island_auto_axi4in_xing_in_aw_mem_2_id),
    .auto_axi4in_xing_in_aw_mem_2_addr(island_auto_axi4in_xing_in_aw_mem_2_addr),
    .auto_axi4in_xing_in_aw_mem_2_len(island_auto_axi4in_xing_in_aw_mem_2_len),
    .auto_axi4in_xing_in_aw_mem_2_size(island_auto_axi4in_xing_in_aw_mem_2_size),
    .auto_axi4in_xing_in_aw_mem_2_burst(island_auto_axi4in_xing_in_aw_mem_2_burst),
    .auto_axi4in_xing_in_aw_mem_2_lock(island_auto_axi4in_xing_in_aw_mem_2_lock),
    .auto_axi4in_xing_in_aw_mem_2_cache(island_auto_axi4in_xing_in_aw_mem_2_cache),
    .auto_axi4in_xing_in_aw_mem_2_prot(island_auto_axi4in_xing_in_aw_mem_2_prot),
    .auto_axi4in_xing_in_aw_mem_2_qos(island_auto_axi4in_xing_in_aw_mem_2_qos),
    .auto_axi4in_xing_in_aw_mem_3_id(island_auto_axi4in_xing_in_aw_mem_3_id),
    .auto_axi4in_xing_in_aw_mem_3_addr(island_auto_axi4in_xing_in_aw_mem_3_addr),
    .auto_axi4in_xing_in_aw_mem_3_len(island_auto_axi4in_xing_in_aw_mem_3_len),
    .auto_axi4in_xing_in_aw_mem_3_size(island_auto_axi4in_xing_in_aw_mem_3_size),
    .auto_axi4in_xing_in_aw_mem_3_burst(island_auto_axi4in_xing_in_aw_mem_3_burst),
    .auto_axi4in_xing_in_aw_mem_3_lock(island_auto_axi4in_xing_in_aw_mem_3_lock),
    .auto_axi4in_xing_in_aw_mem_3_cache(island_auto_axi4in_xing_in_aw_mem_3_cache),
    .auto_axi4in_xing_in_aw_mem_3_prot(island_auto_axi4in_xing_in_aw_mem_3_prot),
    .auto_axi4in_xing_in_aw_mem_3_qos(island_auto_axi4in_xing_in_aw_mem_3_qos),
    .auto_axi4in_xing_in_aw_mem_4_id(island_auto_axi4in_xing_in_aw_mem_4_id),
    .auto_axi4in_xing_in_aw_mem_4_addr(island_auto_axi4in_xing_in_aw_mem_4_addr),
    .auto_axi4in_xing_in_aw_mem_4_len(island_auto_axi4in_xing_in_aw_mem_4_len),
    .auto_axi4in_xing_in_aw_mem_4_size(island_auto_axi4in_xing_in_aw_mem_4_size),
    .auto_axi4in_xing_in_aw_mem_4_burst(island_auto_axi4in_xing_in_aw_mem_4_burst),
    .auto_axi4in_xing_in_aw_mem_4_lock(island_auto_axi4in_xing_in_aw_mem_4_lock),
    .auto_axi4in_xing_in_aw_mem_4_cache(island_auto_axi4in_xing_in_aw_mem_4_cache),
    .auto_axi4in_xing_in_aw_mem_4_prot(island_auto_axi4in_xing_in_aw_mem_4_prot),
    .auto_axi4in_xing_in_aw_mem_4_qos(island_auto_axi4in_xing_in_aw_mem_4_qos),
    .auto_axi4in_xing_in_aw_mem_5_id(island_auto_axi4in_xing_in_aw_mem_5_id),
    .auto_axi4in_xing_in_aw_mem_5_addr(island_auto_axi4in_xing_in_aw_mem_5_addr),
    .auto_axi4in_xing_in_aw_mem_5_len(island_auto_axi4in_xing_in_aw_mem_5_len),
    .auto_axi4in_xing_in_aw_mem_5_size(island_auto_axi4in_xing_in_aw_mem_5_size),
    .auto_axi4in_xing_in_aw_mem_5_burst(island_auto_axi4in_xing_in_aw_mem_5_burst),
    .auto_axi4in_xing_in_aw_mem_5_lock(island_auto_axi4in_xing_in_aw_mem_5_lock),
    .auto_axi4in_xing_in_aw_mem_5_cache(island_auto_axi4in_xing_in_aw_mem_5_cache),
    .auto_axi4in_xing_in_aw_mem_5_prot(island_auto_axi4in_xing_in_aw_mem_5_prot),
    .auto_axi4in_xing_in_aw_mem_5_qos(island_auto_axi4in_xing_in_aw_mem_5_qos),
    .auto_axi4in_xing_in_aw_mem_6_id(island_auto_axi4in_xing_in_aw_mem_6_id),
    .auto_axi4in_xing_in_aw_mem_6_addr(island_auto_axi4in_xing_in_aw_mem_6_addr),
    .auto_axi4in_xing_in_aw_mem_6_len(island_auto_axi4in_xing_in_aw_mem_6_len),
    .auto_axi4in_xing_in_aw_mem_6_size(island_auto_axi4in_xing_in_aw_mem_6_size),
    .auto_axi4in_xing_in_aw_mem_6_burst(island_auto_axi4in_xing_in_aw_mem_6_burst),
    .auto_axi4in_xing_in_aw_mem_6_lock(island_auto_axi4in_xing_in_aw_mem_6_lock),
    .auto_axi4in_xing_in_aw_mem_6_cache(island_auto_axi4in_xing_in_aw_mem_6_cache),
    .auto_axi4in_xing_in_aw_mem_6_prot(island_auto_axi4in_xing_in_aw_mem_6_prot),
    .auto_axi4in_xing_in_aw_mem_6_qos(island_auto_axi4in_xing_in_aw_mem_6_qos),
    .auto_axi4in_xing_in_aw_mem_7_id(island_auto_axi4in_xing_in_aw_mem_7_id),
    .auto_axi4in_xing_in_aw_mem_7_addr(island_auto_axi4in_xing_in_aw_mem_7_addr),
    .auto_axi4in_xing_in_aw_mem_7_len(island_auto_axi4in_xing_in_aw_mem_7_len),
    .auto_axi4in_xing_in_aw_mem_7_size(island_auto_axi4in_xing_in_aw_mem_7_size),
    .auto_axi4in_xing_in_aw_mem_7_burst(island_auto_axi4in_xing_in_aw_mem_7_burst),
    .auto_axi4in_xing_in_aw_mem_7_lock(island_auto_axi4in_xing_in_aw_mem_7_lock),
    .auto_axi4in_xing_in_aw_mem_7_cache(island_auto_axi4in_xing_in_aw_mem_7_cache),
    .auto_axi4in_xing_in_aw_mem_7_prot(island_auto_axi4in_xing_in_aw_mem_7_prot),
    .auto_axi4in_xing_in_aw_mem_7_qos(island_auto_axi4in_xing_in_aw_mem_7_qos),
    .auto_axi4in_xing_in_aw_ridx(island_auto_axi4in_xing_in_aw_ridx),
    .auto_axi4in_xing_in_aw_widx(island_auto_axi4in_xing_in_aw_widx),
    .auto_axi4in_xing_in_aw_safe_ridx_valid(island_auto_axi4in_xing_in_aw_safe_ridx_valid),
    .auto_axi4in_xing_in_aw_safe_widx_valid(island_auto_axi4in_xing_in_aw_safe_widx_valid),
    .auto_axi4in_xing_in_aw_safe_source_reset_n(island_auto_axi4in_xing_in_aw_safe_source_reset_n),
    .auto_axi4in_xing_in_aw_safe_sink_reset_n(island_auto_axi4in_xing_in_aw_safe_sink_reset_n),
    .auto_axi4in_xing_in_w_mem_0_data(island_auto_axi4in_xing_in_w_mem_0_data),
    .auto_axi4in_xing_in_w_mem_0_strb(island_auto_axi4in_xing_in_w_mem_0_strb),
    .auto_axi4in_xing_in_w_mem_0_last(island_auto_axi4in_xing_in_w_mem_0_last),
    .auto_axi4in_xing_in_w_mem_1_data(island_auto_axi4in_xing_in_w_mem_1_data),
    .auto_axi4in_xing_in_w_mem_1_strb(island_auto_axi4in_xing_in_w_mem_1_strb),
    .auto_axi4in_xing_in_w_mem_1_last(island_auto_axi4in_xing_in_w_mem_1_last),
    .auto_axi4in_xing_in_w_mem_2_data(island_auto_axi4in_xing_in_w_mem_2_data),
    .auto_axi4in_xing_in_w_mem_2_strb(island_auto_axi4in_xing_in_w_mem_2_strb),
    .auto_axi4in_xing_in_w_mem_2_last(island_auto_axi4in_xing_in_w_mem_2_last),
    .auto_axi4in_xing_in_w_mem_3_data(island_auto_axi4in_xing_in_w_mem_3_data),
    .auto_axi4in_xing_in_w_mem_3_strb(island_auto_axi4in_xing_in_w_mem_3_strb),
    .auto_axi4in_xing_in_w_mem_3_last(island_auto_axi4in_xing_in_w_mem_3_last),
    .auto_axi4in_xing_in_w_mem_4_data(island_auto_axi4in_xing_in_w_mem_4_data),
    .auto_axi4in_xing_in_w_mem_4_strb(island_auto_axi4in_xing_in_w_mem_4_strb),
    .auto_axi4in_xing_in_w_mem_4_last(island_auto_axi4in_xing_in_w_mem_4_last),
    .auto_axi4in_xing_in_w_mem_5_data(island_auto_axi4in_xing_in_w_mem_5_data),
    .auto_axi4in_xing_in_w_mem_5_strb(island_auto_axi4in_xing_in_w_mem_5_strb),
    .auto_axi4in_xing_in_w_mem_5_last(island_auto_axi4in_xing_in_w_mem_5_last),
    .auto_axi4in_xing_in_w_mem_6_data(island_auto_axi4in_xing_in_w_mem_6_data),
    .auto_axi4in_xing_in_w_mem_6_strb(island_auto_axi4in_xing_in_w_mem_6_strb),
    .auto_axi4in_xing_in_w_mem_6_last(island_auto_axi4in_xing_in_w_mem_6_last),
    .auto_axi4in_xing_in_w_mem_7_data(island_auto_axi4in_xing_in_w_mem_7_data),
    .auto_axi4in_xing_in_w_mem_7_strb(island_auto_axi4in_xing_in_w_mem_7_strb),
    .auto_axi4in_xing_in_w_mem_7_last(island_auto_axi4in_xing_in_w_mem_7_last),
    .auto_axi4in_xing_in_w_ridx(island_auto_axi4in_xing_in_w_ridx),
    .auto_axi4in_xing_in_w_widx(island_auto_axi4in_xing_in_w_widx),
    .auto_axi4in_xing_in_w_safe_ridx_valid(island_auto_axi4in_xing_in_w_safe_ridx_valid),
    .auto_axi4in_xing_in_w_safe_widx_valid(island_auto_axi4in_xing_in_w_safe_widx_valid),
    .auto_axi4in_xing_in_w_safe_source_reset_n(island_auto_axi4in_xing_in_w_safe_source_reset_n),
    .auto_axi4in_xing_in_w_safe_sink_reset_n(island_auto_axi4in_xing_in_w_safe_sink_reset_n),
    .auto_axi4in_xing_in_b_mem_0_id(island_auto_axi4in_xing_in_b_mem_0_id),
    .auto_axi4in_xing_in_b_mem_0_resp(island_auto_axi4in_xing_in_b_mem_0_resp),
    .auto_axi4in_xing_in_b_mem_1_id(island_auto_axi4in_xing_in_b_mem_1_id),
    .auto_axi4in_xing_in_b_mem_1_resp(island_auto_axi4in_xing_in_b_mem_1_resp),
    .auto_axi4in_xing_in_b_mem_2_id(island_auto_axi4in_xing_in_b_mem_2_id),
    .auto_axi4in_xing_in_b_mem_2_resp(island_auto_axi4in_xing_in_b_mem_2_resp),
    .auto_axi4in_xing_in_b_mem_3_id(island_auto_axi4in_xing_in_b_mem_3_id),
    .auto_axi4in_xing_in_b_mem_3_resp(island_auto_axi4in_xing_in_b_mem_3_resp),
    .auto_axi4in_xing_in_b_mem_4_id(island_auto_axi4in_xing_in_b_mem_4_id),
    .auto_axi4in_xing_in_b_mem_4_resp(island_auto_axi4in_xing_in_b_mem_4_resp),
    .auto_axi4in_xing_in_b_mem_5_id(island_auto_axi4in_xing_in_b_mem_5_id),
    .auto_axi4in_xing_in_b_mem_5_resp(island_auto_axi4in_xing_in_b_mem_5_resp),
    .auto_axi4in_xing_in_b_mem_6_id(island_auto_axi4in_xing_in_b_mem_6_id),
    .auto_axi4in_xing_in_b_mem_6_resp(island_auto_axi4in_xing_in_b_mem_6_resp),
    .auto_axi4in_xing_in_b_mem_7_id(island_auto_axi4in_xing_in_b_mem_7_id),
    .auto_axi4in_xing_in_b_mem_7_resp(island_auto_axi4in_xing_in_b_mem_7_resp),
    .auto_axi4in_xing_in_b_ridx(island_auto_axi4in_xing_in_b_ridx),
    .auto_axi4in_xing_in_b_widx(island_auto_axi4in_xing_in_b_widx),
    .auto_axi4in_xing_in_b_safe_ridx_valid(island_auto_axi4in_xing_in_b_safe_ridx_valid),
    .auto_axi4in_xing_in_b_safe_widx_valid(island_auto_axi4in_xing_in_b_safe_widx_valid),
    .auto_axi4in_xing_in_b_safe_source_reset_n(island_auto_axi4in_xing_in_b_safe_source_reset_n),
    .auto_axi4in_xing_in_b_safe_sink_reset_n(island_auto_axi4in_xing_in_b_safe_sink_reset_n),
    .auto_axi4in_xing_in_ar_mem_0_id(island_auto_axi4in_xing_in_ar_mem_0_id),
    .auto_axi4in_xing_in_ar_mem_0_addr(island_auto_axi4in_xing_in_ar_mem_0_addr),
    .auto_axi4in_xing_in_ar_mem_0_len(island_auto_axi4in_xing_in_ar_mem_0_len),
    .auto_axi4in_xing_in_ar_mem_0_size(island_auto_axi4in_xing_in_ar_mem_0_size),
    .auto_axi4in_xing_in_ar_mem_0_burst(island_auto_axi4in_xing_in_ar_mem_0_burst),
    .auto_axi4in_xing_in_ar_mem_0_lock(island_auto_axi4in_xing_in_ar_mem_0_lock),
    .auto_axi4in_xing_in_ar_mem_0_cache(island_auto_axi4in_xing_in_ar_mem_0_cache),
    .auto_axi4in_xing_in_ar_mem_0_prot(island_auto_axi4in_xing_in_ar_mem_0_prot),
    .auto_axi4in_xing_in_ar_mem_0_qos(island_auto_axi4in_xing_in_ar_mem_0_qos),
    .auto_axi4in_xing_in_ar_mem_1_id(island_auto_axi4in_xing_in_ar_mem_1_id),
    .auto_axi4in_xing_in_ar_mem_1_addr(island_auto_axi4in_xing_in_ar_mem_1_addr),
    .auto_axi4in_xing_in_ar_mem_1_len(island_auto_axi4in_xing_in_ar_mem_1_len),
    .auto_axi4in_xing_in_ar_mem_1_size(island_auto_axi4in_xing_in_ar_mem_1_size),
    .auto_axi4in_xing_in_ar_mem_1_burst(island_auto_axi4in_xing_in_ar_mem_1_burst),
    .auto_axi4in_xing_in_ar_mem_1_lock(island_auto_axi4in_xing_in_ar_mem_1_lock),
    .auto_axi4in_xing_in_ar_mem_1_cache(island_auto_axi4in_xing_in_ar_mem_1_cache),
    .auto_axi4in_xing_in_ar_mem_1_prot(island_auto_axi4in_xing_in_ar_mem_1_prot),
    .auto_axi4in_xing_in_ar_mem_1_qos(island_auto_axi4in_xing_in_ar_mem_1_qos),
    .auto_axi4in_xing_in_ar_mem_2_id(island_auto_axi4in_xing_in_ar_mem_2_id),
    .auto_axi4in_xing_in_ar_mem_2_addr(island_auto_axi4in_xing_in_ar_mem_2_addr),
    .auto_axi4in_xing_in_ar_mem_2_len(island_auto_axi4in_xing_in_ar_mem_2_len),
    .auto_axi4in_xing_in_ar_mem_2_size(island_auto_axi4in_xing_in_ar_mem_2_size),
    .auto_axi4in_xing_in_ar_mem_2_burst(island_auto_axi4in_xing_in_ar_mem_2_burst),
    .auto_axi4in_xing_in_ar_mem_2_lock(island_auto_axi4in_xing_in_ar_mem_2_lock),
    .auto_axi4in_xing_in_ar_mem_2_cache(island_auto_axi4in_xing_in_ar_mem_2_cache),
    .auto_axi4in_xing_in_ar_mem_2_prot(island_auto_axi4in_xing_in_ar_mem_2_prot),
    .auto_axi4in_xing_in_ar_mem_2_qos(island_auto_axi4in_xing_in_ar_mem_2_qos),
    .auto_axi4in_xing_in_ar_mem_3_id(island_auto_axi4in_xing_in_ar_mem_3_id),
    .auto_axi4in_xing_in_ar_mem_3_addr(island_auto_axi4in_xing_in_ar_mem_3_addr),
    .auto_axi4in_xing_in_ar_mem_3_len(island_auto_axi4in_xing_in_ar_mem_3_len),
    .auto_axi4in_xing_in_ar_mem_3_size(island_auto_axi4in_xing_in_ar_mem_3_size),
    .auto_axi4in_xing_in_ar_mem_3_burst(island_auto_axi4in_xing_in_ar_mem_3_burst),
    .auto_axi4in_xing_in_ar_mem_3_lock(island_auto_axi4in_xing_in_ar_mem_3_lock),
    .auto_axi4in_xing_in_ar_mem_3_cache(island_auto_axi4in_xing_in_ar_mem_3_cache),
    .auto_axi4in_xing_in_ar_mem_3_prot(island_auto_axi4in_xing_in_ar_mem_3_prot),
    .auto_axi4in_xing_in_ar_mem_3_qos(island_auto_axi4in_xing_in_ar_mem_3_qos),
    .auto_axi4in_xing_in_ar_mem_4_id(island_auto_axi4in_xing_in_ar_mem_4_id),
    .auto_axi4in_xing_in_ar_mem_4_addr(island_auto_axi4in_xing_in_ar_mem_4_addr),
    .auto_axi4in_xing_in_ar_mem_4_len(island_auto_axi4in_xing_in_ar_mem_4_len),
    .auto_axi4in_xing_in_ar_mem_4_size(island_auto_axi4in_xing_in_ar_mem_4_size),
    .auto_axi4in_xing_in_ar_mem_4_burst(island_auto_axi4in_xing_in_ar_mem_4_burst),
    .auto_axi4in_xing_in_ar_mem_4_lock(island_auto_axi4in_xing_in_ar_mem_4_lock),
    .auto_axi4in_xing_in_ar_mem_4_cache(island_auto_axi4in_xing_in_ar_mem_4_cache),
    .auto_axi4in_xing_in_ar_mem_4_prot(island_auto_axi4in_xing_in_ar_mem_4_prot),
    .auto_axi4in_xing_in_ar_mem_4_qos(island_auto_axi4in_xing_in_ar_mem_4_qos),
    .auto_axi4in_xing_in_ar_mem_5_id(island_auto_axi4in_xing_in_ar_mem_5_id),
    .auto_axi4in_xing_in_ar_mem_5_addr(island_auto_axi4in_xing_in_ar_mem_5_addr),
    .auto_axi4in_xing_in_ar_mem_5_len(island_auto_axi4in_xing_in_ar_mem_5_len),
    .auto_axi4in_xing_in_ar_mem_5_size(island_auto_axi4in_xing_in_ar_mem_5_size),
    .auto_axi4in_xing_in_ar_mem_5_burst(island_auto_axi4in_xing_in_ar_mem_5_burst),
    .auto_axi4in_xing_in_ar_mem_5_lock(island_auto_axi4in_xing_in_ar_mem_5_lock),
    .auto_axi4in_xing_in_ar_mem_5_cache(island_auto_axi4in_xing_in_ar_mem_5_cache),
    .auto_axi4in_xing_in_ar_mem_5_prot(island_auto_axi4in_xing_in_ar_mem_5_prot),
    .auto_axi4in_xing_in_ar_mem_5_qos(island_auto_axi4in_xing_in_ar_mem_5_qos),
    .auto_axi4in_xing_in_ar_mem_6_id(island_auto_axi4in_xing_in_ar_mem_6_id),
    .auto_axi4in_xing_in_ar_mem_6_addr(island_auto_axi4in_xing_in_ar_mem_6_addr),
    .auto_axi4in_xing_in_ar_mem_6_len(island_auto_axi4in_xing_in_ar_mem_6_len),
    .auto_axi4in_xing_in_ar_mem_6_size(island_auto_axi4in_xing_in_ar_mem_6_size),
    .auto_axi4in_xing_in_ar_mem_6_burst(island_auto_axi4in_xing_in_ar_mem_6_burst),
    .auto_axi4in_xing_in_ar_mem_6_lock(island_auto_axi4in_xing_in_ar_mem_6_lock),
    .auto_axi4in_xing_in_ar_mem_6_cache(island_auto_axi4in_xing_in_ar_mem_6_cache),
    .auto_axi4in_xing_in_ar_mem_6_prot(island_auto_axi4in_xing_in_ar_mem_6_prot),
    .auto_axi4in_xing_in_ar_mem_6_qos(island_auto_axi4in_xing_in_ar_mem_6_qos),
    .auto_axi4in_xing_in_ar_mem_7_id(island_auto_axi4in_xing_in_ar_mem_7_id),
    .auto_axi4in_xing_in_ar_mem_7_addr(island_auto_axi4in_xing_in_ar_mem_7_addr),
    .auto_axi4in_xing_in_ar_mem_7_len(island_auto_axi4in_xing_in_ar_mem_7_len),
    .auto_axi4in_xing_in_ar_mem_7_size(island_auto_axi4in_xing_in_ar_mem_7_size),
    .auto_axi4in_xing_in_ar_mem_7_burst(island_auto_axi4in_xing_in_ar_mem_7_burst),
    .auto_axi4in_xing_in_ar_mem_7_lock(island_auto_axi4in_xing_in_ar_mem_7_lock),
    .auto_axi4in_xing_in_ar_mem_7_cache(island_auto_axi4in_xing_in_ar_mem_7_cache),
    .auto_axi4in_xing_in_ar_mem_7_prot(island_auto_axi4in_xing_in_ar_mem_7_prot),
    .auto_axi4in_xing_in_ar_mem_7_qos(island_auto_axi4in_xing_in_ar_mem_7_qos),
    .auto_axi4in_xing_in_ar_ridx(island_auto_axi4in_xing_in_ar_ridx),
    .auto_axi4in_xing_in_ar_widx(island_auto_axi4in_xing_in_ar_widx),
    .auto_axi4in_xing_in_ar_safe_ridx_valid(island_auto_axi4in_xing_in_ar_safe_ridx_valid),
    .auto_axi4in_xing_in_ar_safe_widx_valid(island_auto_axi4in_xing_in_ar_safe_widx_valid),
    .auto_axi4in_xing_in_ar_safe_source_reset_n(island_auto_axi4in_xing_in_ar_safe_source_reset_n),
    .auto_axi4in_xing_in_ar_safe_sink_reset_n(island_auto_axi4in_xing_in_ar_safe_sink_reset_n),
    .auto_axi4in_xing_in_r_mem_0_id(island_auto_axi4in_xing_in_r_mem_0_id),
    .auto_axi4in_xing_in_r_mem_0_data(island_auto_axi4in_xing_in_r_mem_0_data),
    .auto_axi4in_xing_in_r_mem_0_resp(island_auto_axi4in_xing_in_r_mem_0_resp),
    .auto_axi4in_xing_in_r_mem_0_last(island_auto_axi4in_xing_in_r_mem_0_last),
    .auto_axi4in_xing_in_r_mem_1_id(island_auto_axi4in_xing_in_r_mem_1_id),
    .auto_axi4in_xing_in_r_mem_1_data(island_auto_axi4in_xing_in_r_mem_1_data),
    .auto_axi4in_xing_in_r_mem_1_resp(island_auto_axi4in_xing_in_r_mem_1_resp),
    .auto_axi4in_xing_in_r_mem_1_last(island_auto_axi4in_xing_in_r_mem_1_last),
    .auto_axi4in_xing_in_r_mem_2_id(island_auto_axi4in_xing_in_r_mem_2_id),
    .auto_axi4in_xing_in_r_mem_2_data(island_auto_axi4in_xing_in_r_mem_2_data),
    .auto_axi4in_xing_in_r_mem_2_resp(island_auto_axi4in_xing_in_r_mem_2_resp),
    .auto_axi4in_xing_in_r_mem_2_last(island_auto_axi4in_xing_in_r_mem_2_last),
    .auto_axi4in_xing_in_r_mem_3_id(island_auto_axi4in_xing_in_r_mem_3_id),
    .auto_axi4in_xing_in_r_mem_3_data(island_auto_axi4in_xing_in_r_mem_3_data),
    .auto_axi4in_xing_in_r_mem_3_resp(island_auto_axi4in_xing_in_r_mem_3_resp),
    .auto_axi4in_xing_in_r_mem_3_last(island_auto_axi4in_xing_in_r_mem_3_last),
    .auto_axi4in_xing_in_r_mem_4_id(island_auto_axi4in_xing_in_r_mem_4_id),
    .auto_axi4in_xing_in_r_mem_4_data(island_auto_axi4in_xing_in_r_mem_4_data),
    .auto_axi4in_xing_in_r_mem_4_resp(island_auto_axi4in_xing_in_r_mem_4_resp),
    .auto_axi4in_xing_in_r_mem_4_last(island_auto_axi4in_xing_in_r_mem_4_last),
    .auto_axi4in_xing_in_r_mem_5_id(island_auto_axi4in_xing_in_r_mem_5_id),
    .auto_axi4in_xing_in_r_mem_5_data(island_auto_axi4in_xing_in_r_mem_5_data),
    .auto_axi4in_xing_in_r_mem_5_resp(island_auto_axi4in_xing_in_r_mem_5_resp),
    .auto_axi4in_xing_in_r_mem_5_last(island_auto_axi4in_xing_in_r_mem_5_last),
    .auto_axi4in_xing_in_r_mem_6_id(island_auto_axi4in_xing_in_r_mem_6_id),
    .auto_axi4in_xing_in_r_mem_6_data(island_auto_axi4in_xing_in_r_mem_6_data),
    .auto_axi4in_xing_in_r_mem_6_resp(island_auto_axi4in_xing_in_r_mem_6_resp),
    .auto_axi4in_xing_in_r_mem_6_last(island_auto_axi4in_xing_in_r_mem_6_last),
    .auto_axi4in_xing_in_r_mem_7_id(island_auto_axi4in_xing_in_r_mem_7_id),
    .auto_axi4in_xing_in_r_mem_7_data(island_auto_axi4in_xing_in_r_mem_7_data),
    .auto_axi4in_xing_in_r_mem_7_resp(island_auto_axi4in_xing_in_r_mem_7_resp),
    .auto_axi4in_xing_in_r_mem_7_last(island_auto_axi4in_xing_in_r_mem_7_last),
    .auto_axi4in_xing_in_r_ridx(island_auto_axi4in_xing_in_r_ridx),
    .auto_axi4in_xing_in_r_widx(island_auto_axi4in_xing_in_r_widx),
    .auto_axi4in_xing_in_r_safe_ridx_valid(island_auto_axi4in_xing_in_r_safe_ridx_valid),
    .auto_axi4in_xing_in_r_safe_widx_valid(island_auto_axi4in_xing_in_r_safe_widx_valid),
    .auto_axi4in_xing_in_r_safe_source_reset_n(island_auto_axi4in_xing_in_r_safe_source_reset_n),
    .auto_axi4in_xing_in_r_safe_sink_reset_n(island_auto_axi4in_xing_in_r_safe_sink_reset_n),
    .io_port_ddr3_addr(island_io_port_ddr3_addr),
    .io_port_ddr3_ba(island_io_port_ddr3_ba),
    .io_port_ddr3_ras_n(island_io_port_ddr3_ras_n),
    .io_port_ddr3_cas_n(island_io_port_ddr3_cas_n),
    .io_port_ddr3_we_n(island_io_port_ddr3_we_n),
    .io_port_ddr3_reset_n(island_io_port_ddr3_reset_n),
    .io_port_ddr3_ck_p(island_io_port_ddr3_ck_p),
    .io_port_ddr3_ck_n(island_io_port_ddr3_ck_n),
    .io_port_ddr3_cke(island_io_port_ddr3_cke),
    .io_port_ddr3_cs_n(island_io_port_ddr3_cs_n),
    .io_port_ddr3_dm(island_io_port_ddr3_dm),
    .io_port_ddr3_odt(island_io_port_ddr3_odt),
    .io_port_ddr3_dq(io_port_ddr3_dq),
    .io_port_ddr3_dqs_n(io_port_ddr3_dqs_n),
    .io_port_ddr3_dqs_p(io_port_ddr3_dqs_p),
    .io_port_sys_clk_i(island_io_port_sys_clk_i),
    .io_port_ui_clk(island_io_port_ui_clk),
    .io_port_ui_clk_sync_rst(island_io_port_ui_clk_sync_rst),
    .io_port_mmcm_locked(island_io_port_mmcm_locked),
    .io_port_aresetn(island_io_port_aresetn),
    .io_port_sys_rst(island_io_port_sys_rst)
  );
  AXI4AsyncCrossingSource axi4asource ( // @[AsyncCrossing.scala 52:33:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310802.4]
    .clock(axi4asource_clock),
    .reset(axi4asource_reset),
    .auto_in_aw_ready(axi4asource_auto_in_aw_ready),
    .auto_in_aw_valid(axi4asource_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4asource_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4asource_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4asource_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4asource_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4asource_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4asource_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4asource_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4asource_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4asource_auto_in_aw_bits_qos),
    .auto_in_w_ready(axi4asource_auto_in_w_ready),
    .auto_in_w_valid(axi4asource_auto_in_w_valid),
    .auto_in_w_bits_data(axi4asource_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4asource_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4asource_auto_in_w_bits_last),
    .auto_in_b_ready(axi4asource_auto_in_b_ready),
    .auto_in_b_valid(axi4asource_auto_in_b_valid),
    .auto_in_b_bits_id(axi4asource_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4asource_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4asource_auto_in_ar_ready),
    .auto_in_ar_valid(axi4asource_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4asource_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4asource_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4asource_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4asource_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4asource_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4asource_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4asource_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4asource_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4asource_auto_in_ar_bits_qos),
    .auto_in_r_ready(axi4asource_auto_in_r_ready),
    .auto_in_r_valid(axi4asource_auto_in_r_valid),
    .auto_in_r_bits_id(axi4asource_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4asource_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4asource_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4asource_auto_in_r_bits_last),
    .auto_out_aw_mem_0_id(axi4asource_auto_out_aw_mem_0_id),
    .auto_out_aw_mem_0_addr(axi4asource_auto_out_aw_mem_0_addr),
    .auto_out_aw_mem_0_len(axi4asource_auto_out_aw_mem_0_len),
    .auto_out_aw_mem_0_size(axi4asource_auto_out_aw_mem_0_size),
    .auto_out_aw_mem_0_burst(axi4asource_auto_out_aw_mem_0_burst),
    .auto_out_aw_mem_0_lock(axi4asource_auto_out_aw_mem_0_lock),
    .auto_out_aw_mem_0_cache(axi4asource_auto_out_aw_mem_0_cache),
    .auto_out_aw_mem_0_prot(axi4asource_auto_out_aw_mem_0_prot),
    .auto_out_aw_mem_0_qos(axi4asource_auto_out_aw_mem_0_qos),
    .auto_out_aw_mem_1_id(axi4asource_auto_out_aw_mem_1_id),
    .auto_out_aw_mem_1_addr(axi4asource_auto_out_aw_mem_1_addr),
    .auto_out_aw_mem_1_len(axi4asource_auto_out_aw_mem_1_len),
    .auto_out_aw_mem_1_size(axi4asource_auto_out_aw_mem_1_size),
    .auto_out_aw_mem_1_burst(axi4asource_auto_out_aw_mem_1_burst),
    .auto_out_aw_mem_1_lock(axi4asource_auto_out_aw_mem_1_lock),
    .auto_out_aw_mem_1_cache(axi4asource_auto_out_aw_mem_1_cache),
    .auto_out_aw_mem_1_prot(axi4asource_auto_out_aw_mem_1_prot),
    .auto_out_aw_mem_1_qos(axi4asource_auto_out_aw_mem_1_qos),
    .auto_out_aw_mem_2_id(axi4asource_auto_out_aw_mem_2_id),
    .auto_out_aw_mem_2_addr(axi4asource_auto_out_aw_mem_2_addr),
    .auto_out_aw_mem_2_len(axi4asource_auto_out_aw_mem_2_len),
    .auto_out_aw_mem_2_size(axi4asource_auto_out_aw_mem_2_size),
    .auto_out_aw_mem_2_burst(axi4asource_auto_out_aw_mem_2_burst),
    .auto_out_aw_mem_2_lock(axi4asource_auto_out_aw_mem_2_lock),
    .auto_out_aw_mem_2_cache(axi4asource_auto_out_aw_mem_2_cache),
    .auto_out_aw_mem_2_prot(axi4asource_auto_out_aw_mem_2_prot),
    .auto_out_aw_mem_2_qos(axi4asource_auto_out_aw_mem_2_qos),
    .auto_out_aw_mem_3_id(axi4asource_auto_out_aw_mem_3_id),
    .auto_out_aw_mem_3_addr(axi4asource_auto_out_aw_mem_3_addr),
    .auto_out_aw_mem_3_len(axi4asource_auto_out_aw_mem_3_len),
    .auto_out_aw_mem_3_size(axi4asource_auto_out_aw_mem_3_size),
    .auto_out_aw_mem_3_burst(axi4asource_auto_out_aw_mem_3_burst),
    .auto_out_aw_mem_3_lock(axi4asource_auto_out_aw_mem_3_lock),
    .auto_out_aw_mem_3_cache(axi4asource_auto_out_aw_mem_3_cache),
    .auto_out_aw_mem_3_prot(axi4asource_auto_out_aw_mem_3_prot),
    .auto_out_aw_mem_3_qos(axi4asource_auto_out_aw_mem_3_qos),
    .auto_out_aw_mem_4_id(axi4asource_auto_out_aw_mem_4_id),
    .auto_out_aw_mem_4_addr(axi4asource_auto_out_aw_mem_4_addr),
    .auto_out_aw_mem_4_len(axi4asource_auto_out_aw_mem_4_len),
    .auto_out_aw_mem_4_size(axi4asource_auto_out_aw_mem_4_size),
    .auto_out_aw_mem_4_burst(axi4asource_auto_out_aw_mem_4_burst),
    .auto_out_aw_mem_4_lock(axi4asource_auto_out_aw_mem_4_lock),
    .auto_out_aw_mem_4_cache(axi4asource_auto_out_aw_mem_4_cache),
    .auto_out_aw_mem_4_prot(axi4asource_auto_out_aw_mem_4_prot),
    .auto_out_aw_mem_4_qos(axi4asource_auto_out_aw_mem_4_qos),
    .auto_out_aw_mem_5_id(axi4asource_auto_out_aw_mem_5_id),
    .auto_out_aw_mem_5_addr(axi4asource_auto_out_aw_mem_5_addr),
    .auto_out_aw_mem_5_len(axi4asource_auto_out_aw_mem_5_len),
    .auto_out_aw_mem_5_size(axi4asource_auto_out_aw_mem_5_size),
    .auto_out_aw_mem_5_burst(axi4asource_auto_out_aw_mem_5_burst),
    .auto_out_aw_mem_5_lock(axi4asource_auto_out_aw_mem_5_lock),
    .auto_out_aw_mem_5_cache(axi4asource_auto_out_aw_mem_5_cache),
    .auto_out_aw_mem_5_prot(axi4asource_auto_out_aw_mem_5_prot),
    .auto_out_aw_mem_5_qos(axi4asource_auto_out_aw_mem_5_qos),
    .auto_out_aw_mem_6_id(axi4asource_auto_out_aw_mem_6_id),
    .auto_out_aw_mem_6_addr(axi4asource_auto_out_aw_mem_6_addr),
    .auto_out_aw_mem_6_len(axi4asource_auto_out_aw_mem_6_len),
    .auto_out_aw_mem_6_size(axi4asource_auto_out_aw_mem_6_size),
    .auto_out_aw_mem_6_burst(axi4asource_auto_out_aw_mem_6_burst),
    .auto_out_aw_mem_6_lock(axi4asource_auto_out_aw_mem_6_lock),
    .auto_out_aw_mem_6_cache(axi4asource_auto_out_aw_mem_6_cache),
    .auto_out_aw_mem_6_prot(axi4asource_auto_out_aw_mem_6_prot),
    .auto_out_aw_mem_6_qos(axi4asource_auto_out_aw_mem_6_qos),
    .auto_out_aw_mem_7_id(axi4asource_auto_out_aw_mem_7_id),
    .auto_out_aw_mem_7_addr(axi4asource_auto_out_aw_mem_7_addr),
    .auto_out_aw_mem_7_len(axi4asource_auto_out_aw_mem_7_len),
    .auto_out_aw_mem_7_size(axi4asource_auto_out_aw_mem_7_size),
    .auto_out_aw_mem_7_burst(axi4asource_auto_out_aw_mem_7_burst),
    .auto_out_aw_mem_7_lock(axi4asource_auto_out_aw_mem_7_lock),
    .auto_out_aw_mem_7_cache(axi4asource_auto_out_aw_mem_7_cache),
    .auto_out_aw_mem_7_prot(axi4asource_auto_out_aw_mem_7_prot),
    .auto_out_aw_mem_7_qos(axi4asource_auto_out_aw_mem_7_qos),
    .auto_out_aw_ridx(axi4asource_auto_out_aw_ridx),
    .auto_out_aw_widx(axi4asource_auto_out_aw_widx),
    .auto_out_aw_safe_ridx_valid(axi4asource_auto_out_aw_safe_ridx_valid),
    .auto_out_aw_safe_widx_valid(axi4asource_auto_out_aw_safe_widx_valid),
    .auto_out_aw_safe_source_reset_n(axi4asource_auto_out_aw_safe_source_reset_n),
    .auto_out_aw_safe_sink_reset_n(axi4asource_auto_out_aw_safe_sink_reset_n),
    .auto_out_w_mem_0_data(axi4asource_auto_out_w_mem_0_data),
    .auto_out_w_mem_0_strb(axi4asource_auto_out_w_mem_0_strb),
    .auto_out_w_mem_0_last(axi4asource_auto_out_w_mem_0_last),
    .auto_out_w_mem_1_data(axi4asource_auto_out_w_mem_1_data),
    .auto_out_w_mem_1_strb(axi4asource_auto_out_w_mem_1_strb),
    .auto_out_w_mem_1_last(axi4asource_auto_out_w_mem_1_last),
    .auto_out_w_mem_2_data(axi4asource_auto_out_w_mem_2_data),
    .auto_out_w_mem_2_strb(axi4asource_auto_out_w_mem_2_strb),
    .auto_out_w_mem_2_last(axi4asource_auto_out_w_mem_2_last),
    .auto_out_w_mem_3_data(axi4asource_auto_out_w_mem_3_data),
    .auto_out_w_mem_3_strb(axi4asource_auto_out_w_mem_3_strb),
    .auto_out_w_mem_3_last(axi4asource_auto_out_w_mem_3_last),
    .auto_out_w_mem_4_data(axi4asource_auto_out_w_mem_4_data),
    .auto_out_w_mem_4_strb(axi4asource_auto_out_w_mem_4_strb),
    .auto_out_w_mem_4_last(axi4asource_auto_out_w_mem_4_last),
    .auto_out_w_mem_5_data(axi4asource_auto_out_w_mem_5_data),
    .auto_out_w_mem_5_strb(axi4asource_auto_out_w_mem_5_strb),
    .auto_out_w_mem_5_last(axi4asource_auto_out_w_mem_5_last),
    .auto_out_w_mem_6_data(axi4asource_auto_out_w_mem_6_data),
    .auto_out_w_mem_6_strb(axi4asource_auto_out_w_mem_6_strb),
    .auto_out_w_mem_6_last(axi4asource_auto_out_w_mem_6_last),
    .auto_out_w_mem_7_data(axi4asource_auto_out_w_mem_7_data),
    .auto_out_w_mem_7_strb(axi4asource_auto_out_w_mem_7_strb),
    .auto_out_w_mem_7_last(axi4asource_auto_out_w_mem_7_last),
    .auto_out_w_ridx(axi4asource_auto_out_w_ridx),
    .auto_out_w_widx(axi4asource_auto_out_w_widx),
    .auto_out_w_safe_ridx_valid(axi4asource_auto_out_w_safe_ridx_valid),
    .auto_out_w_safe_widx_valid(axi4asource_auto_out_w_safe_widx_valid),
    .auto_out_w_safe_source_reset_n(axi4asource_auto_out_w_safe_source_reset_n),
    .auto_out_w_safe_sink_reset_n(axi4asource_auto_out_w_safe_sink_reset_n),
    .auto_out_b_mem_0_id(axi4asource_auto_out_b_mem_0_id),
    .auto_out_b_mem_0_resp(axi4asource_auto_out_b_mem_0_resp),
    .auto_out_b_mem_1_id(axi4asource_auto_out_b_mem_1_id),
    .auto_out_b_mem_1_resp(axi4asource_auto_out_b_mem_1_resp),
    .auto_out_b_mem_2_id(axi4asource_auto_out_b_mem_2_id),
    .auto_out_b_mem_2_resp(axi4asource_auto_out_b_mem_2_resp),
    .auto_out_b_mem_3_id(axi4asource_auto_out_b_mem_3_id),
    .auto_out_b_mem_3_resp(axi4asource_auto_out_b_mem_3_resp),
    .auto_out_b_mem_4_id(axi4asource_auto_out_b_mem_4_id),
    .auto_out_b_mem_4_resp(axi4asource_auto_out_b_mem_4_resp),
    .auto_out_b_mem_5_id(axi4asource_auto_out_b_mem_5_id),
    .auto_out_b_mem_5_resp(axi4asource_auto_out_b_mem_5_resp),
    .auto_out_b_mem_6_id(axi4asource_auto_out_b_mem_6_id),
    .auto_out_b_mem_6_resp(axi4asource_auto_out_b_mem_6_resp),
    .auto_out_b_mem_7_id(axi4asource_auto_out_b_mem_7_id),
    .auto_out_b_mem_7_resp(axi4asource_auto_out_b_mem_7_resp),
    .auto_out_b_ridx(axi4asource_auto_out_b_ridx),
    .auto_out_b_widx(axi4asource_auto_out_b_widx),
    .auto_out_b_safe_ridx_valid(axi4asource_auto_out_b_safe_ridx_valid),
    .auto_out_b_safe_widx_valid(axi4asource_auto_out_b_safe_widx_valid),
    .auto_out_b_safe_source_reset_n(axi4asource_auto_out_b_safe_source_reset_n),
    .auto_out_b_safe_sink_reset_n(axi4asource_auto_out_b_safe_sink_reset_n),
    .auto_out_ar_mem_0_id(axi4asource_auto_out_ar_mem_0_id),
    .auto_out_ar_mem_0_addr(axi4asource_auto_out_ar_mem_0_addr),
    .auto_out_ar_mem_0_len(axi4asource_auto_out_ar_mem_0_len),
    .auto_out_ar_mem_0_size(axi4asource_auto_out_ar_mem_0_size),
    .auto_out_ar_mem_0_burst(axi4asource_auto_out_ar_mem_0_burst),
    .auto_out_ar_mem_0_lock(axi4asource_auto_out_ar_mem_0_lock),
    .auto_out_ar_mem_0_cache(axi4asource_auto_out_ar_mem_0_cache),
    .auto_out_ar_mem_0_prot(axi4asource_auto_out_ar_mem_0_prot),
    .auto_out_ar_mem_0_qos(axi4asource_auto_out_ar_mem_0_qos),
    .auto_out_ar_mem_1_id(axi4asource_auto_out_ar_mem_1_id),
    .auto_out_ar_mem_1_addr(axi4asource_auto_out_ar_mem_1_addr),
    .auto_out_ar_mem_1_len(axi4asource_auto_out_ar_mem_1_len),
    .auto_out_ar_mem_1_size(axi4asource_auto_out_ar_mem_1_size),
    .auto_out_ar_mem_1_burst(axi4asource_auto_out_ar_mem_1_burst),
    .auto_out_ar_mem_1_lock(axi4asource_auto_out_ar_mem_1_lock),
    .auto_out_ar_mem_1_cache(axi4asource_auto_out_ar_mem_1_cache),
    .auto_out_ar_mem_1_prot(axi4asource_auto_out_ar_mem_1_prot),
    .auto_out_ar_mem_1_qos(axi4asource_auto_out_ar_mem_1_qos),
    .auto_out_ar_mem_2_id(axi4asource_auto_out_ar_mem_2_id),
    .auto_out_ar_mem_2_addr(axi4asource_auto_out_ar_mem_2_addr),
    .auto_out_ar_mem_2_len(axi4asource_auto_out_ar_mem_2_len),
    .auto_out_ar_mem_2_size(axi4asource_auto_out_ar_mem_2_size),
    .auto_out_ar_mem_2_burst(axi4asource_auto_out_ar_mem_2_burst),
    .auto_out_ar_mem_2_lock(axi4asource_auto_out_ar_mem_2_lock),
    .auto_out_ar_mem_2_cache(axi4asource_auto_out_ar_mem_2_cache),
    .auto_out_ar_mem_2_prot(axi4asource_auto_out_ar_mem_2_prot),
    .auto_out_ar_mem_2_qos(axi4asource_auto_out_ar_mem_2_qos),
    .auto_out_ar_mem_3_id(axi4asource_auto_out_ar_mem_3_id),
    .auto_out_ar_mem_3_addr(axi4asource_auto_out_ar_mem_3_addr),
    .auto_out_ar_mem_3_len(axi4asource_auto_out_ar_mem_3_len),
    .auto_out_ar_mem_3_size(axi4asource_auto_out_ar_mem_3_size),
    .auto_out_ar_mem_3_burst(axi4asource_auto_out_ar_mem_3_burst),
    .auto_out_ar_mem_3_lock(axi4asource_auto_out_ar_mem_3_lock),
    .auto_out_ar_mem_3_cache(axi4asource_auto_out_ar_mem_3_cache),
    .auto_out_ar_mem_3_prot(axi4asource_auto_out_ar_mem_3_prot),
    .auto_out_ar_mem_3_qos(axi4asource_auto_out_ar_mem_3_qos),
    .auto_out_ar_mem_4_id(axi4asource_auto_out_ar_mem_4_id),
    .auto_out_ar_mem_4_addr(axi4asource_auto_out_ar_mem_4_addr),
    .auto_out_ar_mem_4_len(axi4asource_auto_out_ar_mem_4_len),
    .auto_out_ar_mem_4_size(axi4asource_auto_out_ar_mem_4_size),
    .auto_out_ar_mem_4_burst(axi4asource_auto_out_ar_mem_4_burst),
    .auto_out_ar_mem_4_lock(axi4asource_auto_out_ar_mem_4_lock),
    .auto_out_ar_mem_4_cache(axi4asource_auto_out_ar_mem_4_cache),
    .auto_out_ar_mem_4_prot(axi4asource_auto_out_ar_mem_4_prot),
    .auto_out_ar_mem_4_qos(axi4asource_auto_out_ar_mem_4_qos),
    .auto_out_ar_mem_5_id(axi4asource_auto_out_ar_mem_5_id),
    .auto_out_ar_mem_5_addr(axi4asource_auto_out_ar_mem_5_addr),
    .auto_out_ar_mem_5_len(axi4asource_auto_out_ar_mem_5_len),
    .auto_out_ar_mem_5_size(axi4asource_auto_out_ar_mem_5_size),
    .auto_out_ar_mem_5_burst(axi4asource_auto_out_ar_mem_5_burst),
    .auto_out_ar_mem_5_lock(axi4asource_auto_out_ar_mem_5_lock),
    .auto_out_ar_mem_5_cache(axi4asource_auto_out_ar_mem_5_cache),
    .auto_out_ar_mem_5_prot(axi4asource_auto_out_ar_mem_5_prot),
    .auto_out_ar_mem_5_qos(axi4asource_auto_out_ar_mem_5_qos),
    .auto_out_ar_mem_6_id(axi4asource_auto_out_ar_mem_6_id),
    .auto_out_ar_mem_6_addr(axi4asource_auto_out_ar_mem_6_addr),
    .auto_out_ar_mem_6_len(axi4asource_auto_out_ar_mem_6_len),
    .auto_out_ar_mem_6_size(axi4asource_auto_out_ar_mem_6_size),
    .auto_out_ar_mem_6_burst(axi4asource_auto_out_ar_mem_6_burst),
    .auto_out_ar_mem_6_lock(axi4asource_auto_out_ar_mem_6_lock),
    .auto_out_ar_mem_6_cache(axi4asource_auto_out_ar_mem_6_cache),
    .auto_out_ar_mem_6_prot(axi4asource_auto_out_ar_mem_6_prot),
    .auto_out_ar_mem_6_qos(axi4asource_auto_out_ar_mem_6_qos),
    .auto_out_ar_mem_7_id(axi4asource_auto_out_ar_mem_7_id),
    .auto_out_ar_mem_7_addr(axi4asource_auto_out_ar_mem_7_addr),
    .auto_out_ar_mem_7_len(axi4asource_auto_out_ar_mem_7_len),
    .auto_out_ar_mem_7_size(axi4asource_auto_out_ar_mem_7_size),
    .auto_out_ar_mem_7_burst(axi4asource_auto_out_ar_mem_7_burst),
    .auto_out_ar_mem_7_lock(axi4asource_auto_out_ar_mem_7_lock),
    .auto_out_ar_mem_7_cache(axi4asource_auto_out_ar_mem_7_cache),
    .auto_out_ar_mem_7_prot(axi4asource_auto_out_ar_mem_7_prot),
    .auto_out_ar_mem_7_qos(axi4asource_auto_out_ar_mem_7_qos),
    .auto_out_ar_ridx(axi4asource_auto_out_ar_ridx),
    .auto_out_ar_widx(axi4asource_auto_out_ar_widx),
    .auto_out_ar_safe_ridx_valid(axi4asource_auto_out_ar_safe_ridx_valid),
    .auto_out_ar_safe_widx_valid(axi4asource_auto_out_ar_safe_widx_valid),
    .auto_out_ar_safe_source_reset_n(axi4asource_auto_out_ar_safe_source_reset_n),
    .auto_out_ar_safe_sink_reset_n(axi4asource_auto_out_ar_safe_sink_reset_n),
    .auto_out_r_mem_0_id(axi4asource_auto_out_r_mem_0_id),
    .auto_out_r_mem_0_data(axi4asource_auto_out_r_mem_0_data),
    .auto_out_r_mem_0_resp(axi4asource_auto_out_r_mem_0_resp),
    .auto_out_r_mem_0_last(axi4asource_auto_out_r_mem_0_last),
    .auto_out_r_mem_1_id(axi4asource_auto_out_r_mem_1_id),
    .auto_out_r_mem_1_data(axi4asource_auto_out_r_mem_1_data),
    .auto_out_r_mem_1_resp(axi4asource_auto_out_r_mem_1_resp),
    .auto_out_r_mem_1_last(axi4asource_auto_out_r_mem_1_last),
    .auto_out_r_mem_2_id(axi4asource_auto_out_r_mem_2_id),
    .auto_out_r_mem_2_data(axi4asource_auto_out_r_mem_2_data),
    .auto_out_r_mem_2_resp(axi4asource_auto_out_r_mem_2_resp),
    .auto_out_r_mem_2_last(axi4asource_auto_out_r_mem_2_last),
    .auto_out_r_mem_3_id(axi4asource_auto_out_r_mem_3_id),
    .auto_out_r_mem_3_data(axi4asource_auto_out_r_mem_3_data),
    .auto_out_r_mem_3_resp(axi4asource_auto_out_r_mem_3_resp),
    .auto_out_r_mem_3_last(axi4asource_auto_out_r_mem_3_last),
    .auto_out_r_mem_4_id(axi4asource_auto_out_r_mem_4_id),
    .auto_out_r_mem_4_data(axi4asource_auto_out_r_mem_4_data),
    .auto_out_r_mem_4_resp(axi4asource_auto_out_r_mem_4_resp),
    .auto_out_r_mem_4_last(axi4asource_auto_out_r_mem_4_last),
    .auto_out_r_mem_5_id(axi4asource_auto_out_r_mem_5_id),
    .auto_out_r_mem_5_data(axi4asource_auto_out_r_mem_5_data),
    .auto_out_r_mem_5_resp(axi4asource_auto_out_r_mem_5_resp),
    .auto_out_r_mem_5_last(axi4asource_auto_out_r_mem_5_last),
    .auto_out_r_mem_6_id(axi4asource_auto_out_r_mem_6_id),
    .auto_out_r_mem_6_data(axi4asource_auto_out_r_mem_6_data),
    .auto_out_r_mem_6_resp(axi4asource_auto_out_r_mem_6_resp),
    .auto_out_r_mem_6_last(axi4asource_auto_out_r_mem_6_last),
    .auto_out_r_mem_7_id(axi4asource_auto_out_r_mem_7_id),
    .auto_out_r_mem_7_data(axi4asource_auto_out_r_mem_7_data),
    .auto_out_r_mem_7_resp(axi4asource_auto_out_r_mem_7_resp),
    .auto_out_r_mem_7_last(axi4asource_auto_out_r_mem_7_last),
    .auto_out_r_ridx(axi4asource_auto_out_r_ridx),
    .auto_out_r_widx(axi4asource_auto_out_r_widx),
    .auto_out_r_safe_ridx_valid(axi4asource_auto_out_r_safe_ridx_valid),
    .auto_out_r_safe_widx_valid(axi4asource_auto_out_r_safe_widx_valid),
    .auto_out_r_safe_source_reset_n(axi4asource_auto_out_r_safe_source_reset_n),
    .auto_out_r_safe_sink_reset_n(axi4asource_auto_out_r_safe_sink_reset_n)
  );
  assign auto_buffer_in_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign auto_buffer_in_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign auto_buffer_in_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign auto_buffer_in_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign auto_buffer_in_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign auto_buffer_in_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign auto_buffer_in_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign auto_buffer_in_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign auto_buffer_in_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign io_port_ddr3_addr = island_io_port_ddr3_addr; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_ba = island_io_port_ddr3_ba; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_ras_n = island_io_port_ddr3_ras_n; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_cas_n = island_io_port_ddr3_cas_n; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_we_n = island_io_port_ddr3_we_n; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_reset_n = island_io_port_ddr3_reset_n; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_ck_p = island_io_port_ddr3_ck_p; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_ck_n = island_io_port_ddr3_ck_n; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_cke = island_io_port_ddr3_cke; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_cs_n = island_io_port_ddr3_cs_n; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_dm = island_io_port_ddr3_dm; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ddr3_odt = island_io_port_ddr3_odt; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ui_clk = island_io_port_ui_clk; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_ui_clk_sync_rst = island_io_port_ui_clk_sync_rst; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign io_port_mmcm_locked = island_io_port_mmcm_locked; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign buffer_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310773.4]
  assign buffer_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310774.4]
  assign buffer_auto_in_a_valid = auto_buffer_in_a_valid; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign buffer_auto_in_a_bits_opcode = auto_buffer_in_a_bits_opcode; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign buffer_auto_in_a_bits_size = auto_buffer_in_a_bits_size; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign buffer_auto_in_a_bits_source = auto_buffer_in_a_bits_source; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign buffer_auto_in_a_bits_address = auto_buffer_in_a_bits_address; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign buffer_auto_in_a_bits_mask = auto_buffer_in_a_bits_mask; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign buffer_auto_in_a_bits_data = auto_buffer_in_a_bits_data; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign buffer_auto_in_d_ready = auto_buffer_in_d_ready; // @[LazyModule.scala 173:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310820.4]
  assign buffer_auto_out_a_ready = toaxi4_auto_in_a_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign buffer_auto_out_d_valid = toaxi4_auto_in_d_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign buffer_auto_out_d_bits_opcode = toaxi4_auto_in_d_bits_opcode; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign buffer_auto_out_d_bits_size = toaxi4_auto_in_d_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign buffer_auto_out_d_bits_source = toaxi4_auto_in_d_bits_source; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign buffer_auto_out_d_bits_denied = toaxi4_auto_in_d_bits_denied; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign buffer_auto_out_d_bits_data = toaxi4_auto_in_d_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign buffer_auto_out_d_bits_corrupt = toaxi4_auto_in_d_bits_corrupt; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310779.4]
  assign toaxi4_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310780.4]
  assign toaxi4_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310813.4]
  assign toaxi4_auto_out_aw_ready = indexer_auto_in_aw_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_w_ready = indexer_auto_in_w_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_b_valid = indexer_auto_in_b_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_b_bits_id = indexer_auto_in_b_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_b_bits_resp = indexer_auto_in_b_bits_resp; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_b_bits_user = indexer_auto_in_b_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_ar_ready = indexer_auto_in_ar_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_r_valid = indexer_auto_in_r_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_r_bits_id = indexer_auto_in_r_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_r_bits_data = indexer_auto_in_r_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_r_bits_resp = indexer_auto_in_r_bits_resp; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_r_bits_user = indexer_auto_in_r_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign toaxi4_auto_out_r_bits_last = indexer_auto_in_r_bits_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_valid = toaxi4_auto_out_aw_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_id = toaxi4_auto_out_aw_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_addr = toaxi4_auto_out_aw_bits_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_len = toaxi4_auto_out_aw_bits_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_size = toaxi4_auto_out_aw_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_burst = toaxi4_auto_out_aw_bits_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_lock = toaxi4_auto_out_aw_bits_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_cache = toaxi4_auto_out_aw_bits_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_prot = toaxi4_auto_out_aw_bits_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_qos = toaxi4_auto_out_aw_bits_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_aw_bits_user = toaxi4_auto_out_aw_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_w_valid = toaxi4_auto_out_w_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_w_bits_data = toaxi4_auto_out_w_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_w_bits_strb = toaxi4_auto_out_w_bits_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_w_bits_last = toaxi4_auto_out_w_bits_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_b_ready = toaxi4_auto_out_b_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_valid = toaxi4_auto_out_ar_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_id = toaxi4_auto_out_ar_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_addr = toaxi4_auto_out_ar_bits_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_len = toaxi4_auto_out_ar_bits_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_size = toaxi4_auto_out_ar_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_burst = toaxi4_auto_out_ar_bits_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_lock = toaxi4_auto_out_ar_bits_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_cache = toaxi4_auto_out_ar_bits_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_prot = toaxi4_auto_out_ar_bits_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_qos = toaxi4_auto_out_ar_bits_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_ar_bits_user = toaxi4_auto_out_ar_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_in_r_ready = toaxi4_auto_out_r_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310814.4]
  assign indexer_auto_out_aw_ready = deint_auto_in_aw_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_w_ready = deint_auto_in_w_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_b_valid = deint_auto_in_b_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_b_bits_id = deint_auto_in_b_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_b_bits_resp = deint_auto_in_b_bits_resp; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_b_bits_user = deint_auto_in_b_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_ar_ready = deint_auto_in_ar_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_r_valid = deint_auto_in_r_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_r_bits_id = deint_auto_in_r_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_r_bits_data = deint_auto_in_r_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_r_bits_resp = deint_auto_in_r_bits_resp; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_r_bits_user = deint_auto_in_r_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign indexer_auto_out_r_bits_last = deint_auto_in_r_bits_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310791.4]
  assign deint_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310792.4]
  assign deint_auto_in_aw_valid = indexer_auto_out_aw_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_id = indexer_auto_out_aw_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_addr = indexer_auto_out_aw_bits_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_len = indexer_auto_out_aw_bits_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_size = indexer_auto_out_aw_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_burst = indexer_auto_out_aw_bits_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_lock = indexer_auto_out_aw_bits_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_cache = indexer_auto_out_aw_bits_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_prot = indexer_auto_out_aw_bits_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_qos = indexer_auto_out_aw_bits_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_aw_bits_user = indexer_auto_out_aw_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_w_valid = indexer_auto_out_w_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_w_bits_data = indexer_auto_out_w_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_w_bits_strb = indexer_auto_out_w_bits_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_w_bits_last = indexer_auto_out_w_bits_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_b_ready = indexer_auto_out_b_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_valid = indexer_auto_out_ar_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_id = indexer_auto_out_ar_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_addr = indexer_auto_out_ar_bits_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_len = indexer_auto_out_ar_bits_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_size = indexer_auto_out_ar_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_burst = indexer_auto_out_ar_bits_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_lock = indexer_auto_out_ar_bits_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_cache = indexer_auto_out_ar_bits_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_prot = indexer_auto_out_ar_bits_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_qos = indexer_auto_out_ar_bits_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_ar_bits_user = indexer_auto_out_ar_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_in_r_ready = indexer_auto_out_r_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310815.4]
  assign deint_auto_out_aw_ready = yank_auto_in_aw_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_w_ready = yank_auto_in_w_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_b_valid = yank_auto_in_b_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_b_bits_id = yank_auto_in_b_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_b_bits_resp = yank_auto_in_b_bits_resp; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_b_bits_user = yank_auto_in_b_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_ar_ready = yank_auto_in_ar_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_r_valid = yank_auto_in_r_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_r_bits_id = yank_auto_in_r_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_r_bits_data = yank_auto_in_r_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_r_bits_resp = yank_auto_in_r_bits_resp; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_r_bits_user = yank_auto_in_r_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign deint_auto_out_r_bits_last = yank_auto_in_r_bits_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310797.4]
  assign yank_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310798.4]
  assign yank_auto_in_aw_valid = deint_auto_out_aw_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_id = deint_auto_out_aw_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_addr = deint_auto_out_aw_bits_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_len = deint_auto_out_aw_bits_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_size = deint_auto_out_aw_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_burst = deint_auto_out_aw_bits_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_lock = deint_auto_out_aw_bits_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_cache = deint_auto_out_aw_bits_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_prot = deint_auto_out_aw_bits_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_qos = deint_auto_out_aw_bits_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_aw_bits_user = deint_auto_out_aw_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_w_valid = deint_auto_out_w_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_w_bits_data = deint_auto_out_w_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_w_bits_strb = deint_auto_out_w_bits_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_w_bits_last = deint_auto_out_w_bits_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_b_ready = deint_auto_out_b_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_valid = deint_auto_out_ar_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_id = deint_auto_out_ar_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_addr = deint_auto_out_ar_bits_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_len = deint_auto_out_ar_bits_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_size = deint_auto_out_ar_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_burst = deint_auto_out_ar_bits_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_lock = deint_auto_out_ar_bits_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_cache = deint_auto_out_ar_bits_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_prot = deint_auto_out_ar_bits_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_qos = deint_auto_out_ar_bits_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_ar_bits_user = deint_auto_out_ar_bits_user; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_in_r_ready = deint_auto_out_r_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310816.4]
  assign yank_auto_out_aw_ready = axi4asource_auto_in_aw_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_w_ready = axi4asource_auto_in_w_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_b_valid = axi4asource_auto_in_b_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_b_bits_id = axi4asource_auto_in_b_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_b_bits_resp = axi4asource_auto_in_b_bits_resp; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_ar_ready = axi4asource_auto_in_ar_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_r_valid = axi4asource_auto_in_r_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_r_bits_id = axi4asource_auto_in_r_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_r_bits_data = axi4asource_auto_in_r_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_r_bits_resp = axi4asource_auto_in_r_bits_resp; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign yank_auto_out_r_bits_last = axi4asource_auto_in_r_bits_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_id = axi4asource_auto_out_aw_mem_0_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_addr = axi4asource_auto_out_aw_mem_0_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_len = axi4asource_auto_out_aw_mem_0_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_size = axi4asource_auto_out_aw_mem_0_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_burst = axi4asource_auto_out_aw_mem_0_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_lock = axi4asource_auto_out_aw_mem_0_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_cache = axi4asource_auto_out_aw_mem_0_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_prot = axi4asource_auto_out_aw_mem_0_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_0_qos = axi4asource_auto_out_aw_mem_0_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_id = axi4asource_auto_out_aw_mem_1_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_addr = axi4asource_auto_out_aw_mem_1_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_len = axi4asource_auto_out_aw_mem_1_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_size = axi4asource_auto_out_aw_mem_1_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_burst = axi4asource_auto_out_aw_mem_1_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_lock = axi4asource_auto_out_aw_mem_1_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_cache = axi4asource_auto_out_aw_mem_1_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_prot = axi4asource_auto_out_aw_mem_1_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_1_qos = axi4asource_auto_out_aw_mem_1_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_id = axi4asource_auto_out_aw_mem_2_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_addr = axi4asource_auto_out_aw_mem_2_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_len = axi4asource_auto_out_aw_mem_2_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_size = axi4asource_auto_out_aw_mem_2_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_burst = axi4asource_auto_out_aw_mem_2_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_lock = axi4asource_auto_out_aw_mem_2_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_cache = axi4asource_auto_out_aw_mem_2_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_prot = axi4asource_auto_out_aw_mem_2_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_2_qos = axi4asource_auto_out_aw_mem_2_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_id = axi4asource_auto_out_aw_mem_3_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_addr = axi4asource_auto_out_aw_mem_3_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_len = axi4asource_auto_out_aw_mem_3_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_size = axi4asource_auto_out_aw_mem_3_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_burst = axi4asource_auto_out_aw_mem_3_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_lock = axi4asource_auto_out_aw_mem_3_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_cache = axi4asource_auto_out_aw_mem_3_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_prot = axi4asource_auto_out_aw_mem_3_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_3_qos = axi4asource_auto_out_aw_mem_3_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_id = axi4asource_auto_out_aw_mem_4_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_addr = axi4asource_auto_out_aw_mem_4_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_len = axi4asource_auto_out_aw_mem_4_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_size = axi4asource_auto_out_aw_mem_4_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_burst = axi4asource_auto_out_aw_mem_4_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_lock = axi4asource_auto_out_aw_mem_4_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_cache = axi4asource_auto_out_aw_mem_4_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_prot = axi4asource_auto_out_aw_mem_4_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_4_qos = axi4asource_auto_out_aw_mem_4_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_id = axi4asource_auto_out_aw_mem_5_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_addr = axi4asource_auto_out_aw_mem_5_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_len = axi4asource_auto_out_aw_mem_5_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_size = axi4asource_auto_out_aw_mem_5_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_burst = axi4asource_auto_out_aw_mem_5_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_lock = axi4asource_auto_out_aw_mem_5_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_cache = axi4asource_auto_out_aw_mem_5_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_prot = axi4asource_auto_out_aw_mem_5_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_5_qos = axi4asource_auto_out_aw_mem_5_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_id = axi4asource_auto_out_aw_mem_6_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_addr = axi4asource_auto_out_aw_mem_6_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_len = axi4asource_auto_out_aw_mem_6_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_size = axi4asource_auto_out_aw_mem_6_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_burst = axi4asource_auto_out_aw_mem_6_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_lock = axi4asource_auto_out_aw_mem_6_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_cache = axi4asource_auto_out_aw_mem_6_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_prot = axi4asource_auto_out_aw_mem_6_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_6_qos = axi4asource_auto_out_aw_mem_6_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_id = axi4asource_auto_out_aw_mem_7_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_addr = axi4asource_auto_out_aw_mem_7_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_len = axi4asource_auto_out_aw_mem_7_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_size = axi4asource_auto_out_aw_mem_7_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_burst = axi4asource_auto_out_aw_mem_7_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_lock = axi4asource_auto_out_aw_mem_7_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_cache = axi4asource_auto_out_aw_mem_7_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_prot = axi4asource_auto_out_aw_mem_7_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_mem_7_qos = axi4asource_auto_out_aw_mem_7_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_widx = axi4asource_auto_out_aw_widx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_safe_widx_valid = axi4asource_auto_out_aw_safe_widx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_aw_safe_source_reset_n = axi4asource_auto_out_aw_safe_source_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_0_data = axi4asource_auto_out_w_mem_0_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_0_strb = axi4asource_auto_out_w_mem_0_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_0_last = axi4asource_auto_out_w_mem_0_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_1_data = axi4asource_auto_out_w_mem_1_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_1_strb = axi4asource_auto_out_w_mem_1_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_1_last = axi4asource_auto_out_w_mem_1_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_2_data = axi4asource_auto_out_w_mem_2_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_2_strb = axi4asource_auto_out_w_mem_2_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_2_last = axi4asource_auto_out_w_mem_2_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_3_data = axi4asource_auto_out_w_mem_3_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_3_strb = axi4asource_auto_out_w_mem_3_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_3_last = axi4asource_auto_out_w_mem_3_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_4_data = axi4asource_auto_out_w_mem_4_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_4_strb = axi4asource_auto_out_w_mem_4_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_4_last = axi4asource_auto_out_w_mem_4_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_5_data = axi4asource_auto_out_w_mem_5_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_5_strb = axi4asource_auto_out_w_mem_5_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_5_last = axi4asource_auto_out_w_mem_5_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_6_data = axi4asource_auto_out_w_mem_6_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_6_strb = axi4asource_auto_out_w_mem_6_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_6_last = axi4asource_auto_out_w_mem_6_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_7_data = axi4asource_auto_out_w_mem_7_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_7_strb = axi4asource_auto_out_w_mem_7_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_mem_7_last = axi4asource_auto_out_w_mem_7_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_widx = axi4asource_auto_out_w_widx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_safe_widx_valid = axi4asource_auto_out_w_safe_widx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_w_safe_source_reset_n = axi4asource_auto_out_w_safe_source_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_b_ridx = axi4asource_auto_out_b_ridx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_b_safe_ridx_valid = axi4asource_auto_out_b_safe_ridx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_b_safe_sink_reset_n = axi4asource_auto_out_b_safe_sink_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_id = axi4asource_auto_out_ar_mem_0_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_addr = axi4asource_auto_out_ar_mem_0_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_len = axi4asource_auto_out_ar_mem_0_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_size = axi4asource_auto_out_ar_mem_0_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_burst = axi4asource_auto_out_ar_mem_0_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_lock = axi4asource_auto_out_ar_mem_0_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_cache = axi4asource_auto_out_ar_mem_0_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_prot = axi4asource_auto_out_ar_mem_0_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_0_qos = axi4asource_auto_out_ar_mem_0_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_id = axi4asource_auto_out_ar_mem_1_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_addr = axi4asource_auto_out_ar_mem_1_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_len = axi4asource_auto_out_ar_mem_1_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_size = axi4asource_auto_out_ar_mem_1_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_burst = axi4asource_auto_out_ar_mem_1_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_lock = axi4asource_auto_out_ar_mem_1_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_cache = axi4asource_auto_out_ar_mem_1_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_prot = axi4asource_auto_out_ar_mem_1_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_1_qos = axi4asource_auto_out_ar_mem_1_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_id = axi4asource_auto_out_ar_mem_2_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_addr = axi4asource_auto_out_ar_mem_2_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_len = axi4asource_auto_out_ar_mem_2_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_size = axi4asource_auto_out_ar_mem_2_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_burst = axi4asource_auto_out_ar_mem_2_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_lock = axi4asource_auto_out_ar_mem_2_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_cache = axi4asource_auto_out_ar_mem_2_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_prot = axi4asource_auto_out_ar_mem_2_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_2_qos = axi4asource_auto_out_ar_mem_2_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_id = axi4asource_auto_out_ar_mem_3_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_addr = axi4asource_auto_out_ar_mem_3_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_len = axi4asource_auto_out_ar_mem_3_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_size = axi4asource_auto_out_ar_mem_3_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_burst = axi4asource_auto_out_ar_mem_3_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_lock = axi4asource_auto_out_ar_mem_3_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_cache = axi4asource_auto_out_ar_mem_3_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_prot = axi4asource_auto_out_ar_mem_3_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_3_qos = axi4asource_auto_out_ar_mem_3_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_id = axi4asource_auto_out_ar_mem_4_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_addr = axi4asource_auto_out_ar_mem_4_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_len = axi4asource_auto_out_ar_mem_4_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_size = axi4asource_auto_out_ar_mem_4_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_burst = axi4asource_auto_out_ar_mem_4_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_lock = axi4asource_auto_out_ar_mem_4_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_cache = axi4asource_auto_out_ar_mem_4_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_prot = axi4asource_auto_out_ar_mem_4_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_4_qos = axi4asource_auto_out_ar_mem_4_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_id = axi4asource_auto_out_ar_mem_5_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_addr = axi4asource_auto_out_ar_mem_5_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_len = axi4asource_auto_out_ar_mem_5_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_size = axi4asource_auto_out_ar_mem_5_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_burst = axi4asource_auto_out_ar_mem_5_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_lock = axi4asource_auto_out_ar_mem_5_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_cache = axi4asource_auto_out_ar_mem_5_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_prot = axi4asource_auto_out_ar_mem_5_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_5_qos = axi4asource_auto_out_ar_mem_5_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_id = axi4asource_auto_out_ar_mem_6_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_addr = axi4asource_auto_out_ar_mem_6_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_len = axi4asource_auto_out_ar_mem_6_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_size = axi4asource_auto_out_ar_mem_6_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_burst = axi4asource_auto_out_ar_mem_6_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_lock = axi4asource_auto_out_ar_mem_6_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_cache = axi4asource_auto_out_ar_mem_6_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_prot = axi4asource_auto_out_ar_mem_6_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_6_qos = axi4asource_auto_out_ar_mem_6_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_id = axi4asource_auto_out_ar_mem_7_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_addr = axi4asource_auto_out_ar_mem_7_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_len = axi4asource_auto_out_ar_mem_7_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_size = axi4asource_auto_out_ar_mem_7_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_burst = axi4asource_auto_out_ar_mem_7_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_lock = axi4asource_auto_out_ar_mem_7_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_cache = axi4asource_auto_out_ar_mem_7_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_prot = axi4asource_auto_out_ar_mem_7_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_mem_7_qos = axi4asource_auto_out_ar_mem_7_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_widx = axi4asource_auto_out_ar_widx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_safe_widx_valid = axi4asource_auto_out_ar_safe_widx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_ar_safe_source_reset_n = axi4asource_auto_out_ar_safe_source_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_r_ridx = axi4asource_auto_out_r_ridx; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_r_safe_ridx_valid = axi4asource_auto_out_r_safe_ridx_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_auto_axi4in_xing_in_r_safe_sink_reset_n = axi4asource_auto_out_r_safe_sink_reset_n; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310818.4]
  assign island_io_port_sys_clk_i = io_port_sys_clk_i; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign island_io_port_aresetn = io_port_aresetn; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign island_io_port_sys_rst = io_port_sys_rst; // @[XilinxVC707MIG.scala 168:13:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310821.4]
  assign axi4asource_clock = clock; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310806.4]
  assign axi4asource_reset = reset; // @[:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310807.4]
  assign axi4asource_auto_in_aw_valid = yank_auto_out_aw_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_id = yank_auto_out_aw_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_addr = yank_auto_out_aw_bits_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_len = yank_auto_out_aw_bits_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_size = yank_auto_out_aw_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_burst = yank_auto_out_aw_bits_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_lock = yank_auto_out_aw_bits_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_cache = yank_auto_out_aw_bits_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_prot = yank_auto_out_aw_bits_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_aw_bits_qos = yank_auto_out_aw_bits_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_w_valid = yank_auto_out_w_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_w_bits_data = yank_auto_out_w_bits_data; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_w_bits_strb = yank_auto_out_w_bits_strb; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_w_bits_last = yank_auto_out_w_bits_last; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_b_ready = yank_auto_out_b_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_valid = yank_auto_out_ar_valid; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_id = yank_auto_out_ar_bits_id; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_addr = yank_auto_out_ar_bits_addr; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_len = yank_auto_out_ar_bits_len; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_size = yank_auto_out_ar_bits_size; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_burst = yank_auto_out_ar_bits_burst; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_lock = yank_auto_out_ar_bits_lock; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_cache = yank_auto_out_ar_bits_cache; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_prot = yank_auto_out_ar_bits_prot; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_ar_bits_qos = yank_auto_out_ar_bits_qos; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_in_r_ready = yank_auto_out_r_ready; // @[LazyModule.scala 167:57:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310817.4]
  assign axi4asource_auto_out_aw_ridx = island_auto_axi4in_xing_in_aw_ridx; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_aw_safe_ridx_valid = island_auto_axi4in_xing_in_aw_safe_ridx_valid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_aw_safe_sink_reset_n = island_auto_axi4in_xing_in_aw_safe_sink_reset_n; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_w_ridx = island_auto_axi4in_xing_in_w_ridx; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_w_safe_ridx_valid = island_auto_axi4in_xing_in_w_safe_ridx_valid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_w_safe_sink_reset_n = island_auto_axi4in_xing_in_w_safe_sink_reset_n; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_0_id = island_auto_axi4in_xing_in_b_mem_0_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_0_resp = island_auto_axi4in_xing_in_b_mem_0_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_1_id = island_auto_axi4in_xing_in_b_mem_1_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_1_resp = island_auto_axi4in_xing_in_b_mem_1_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_2_id = island_auto_axi4in_xing_in_b_mem_2_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_2_resp = island_auto_axi4in_xing_in_b_mem_2_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_3_id = island_auto_axi4in_xing_in_b_mem_3_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_3_resp = island_auto_axi4in_xing_in_b_mem_3_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_4_id = island_auto_axi4in_xing_in_b_mem_4_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_4_resp = island_auto_axi4in_xing_in_b_mem_4_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_5_id = island_auto_axi4in_xing_in_b_mem_5_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_5_resp = island_auto_axi4in_xing_in_b_mem_5_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_6_id = island_auto_axi4in_xing_in_b_mem_6_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_6_resp = island_auto_axi4in_xing_in_b_mem_6_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_7_id = island_auto_axi4in_xing_in_b_mem_7_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_mem_7_resp = island_auto_axi4in_xing_in_b_mem_7_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_widx = island_auto_axi4in_xing_in_b_widx; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_safe_widx_valid = island_auto_axi4in_xing_in_b_safe_widx_valid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_b_safe_source_reset_n = island_auto_axi4in_xing_in_b_safe_source_reset_n; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_ar_ridx = island_auto_axi4in_xing_in_ar_ridx; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_ar_safe_ridx_valid = island_auto_axi4in_xing_in_ar_safe_ridx_valid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_ar_safe_sink_reset_n = island_auto_axi4in_xing_in_ar_safe_sink_reset_n; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_0_id = island_auto_axi4in_xing_in_r_mem_0_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_0_data = island_auto_axi4in_xing_in_r_mem_0_data; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_0_resp = island_auto_axi4in_xing_in_r_mem_0_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_0_last = island_auto_axi4in_xing_in_r_mem_0_last; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_1_id = island_auto_axi4in_xing_in_r_mem_1_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_1_data = island_auto_axi4in_xing_in_r_mem_1_data; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_1_resp = island_auto_axi4in_xing_in_r_mem_1_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_1_last = island_auto_axi4in_xing_in_r_mem_1_last; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_2_id = island_auto_axi4in_xing_in_r_mem_2_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_2_data = island_auto_axi4in_xing_in_r_mem_2_data; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_2_resp = island_auto_axi4in_xing_in_r_mem_2_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_2_last = island_auto_axi4in_xing_in_r_mem_2_last; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_3_id = island_auto_axi4in_xing_in_r_mem_3_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_3_data = island_auto_axi4in_xing_in_r_mem_3_data; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_3_resp = island_auto_axi4in_xing_in_r_mem_3_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_3_last = island_auto_axi4in_xing_in_r_mem_3_last; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_4_id = island_auto_axi4in_xing_in_r_mem_4_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_4_data = island_auto_axi4in_xing_in_r_mem_4_data; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_4_resp = island_auto_axi4in_xing_in_r_mem_4_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_4_last = island_auto_axi4in_xing_in_r_mem_4_last; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_5_id = island_auto_axi4in_xing_in_r_mem_5_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_5_data = island_auto_axi4in_xing_in_r_mem_5_data; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_5_resp = island_auto_axi4in_xing_in_r_mem_5_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_5_last = island_auto_axi4in_xing_in_r_mem_5_last; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_6_id = island_auto_axi4in_xing_in_r_mem_6_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_6_data = island_auto_axi4in_xing_in_r_mem_6_data; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_6_resp = island_auto_axi4in_xing_in_r_mem_6_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_6_last = island_auto_axi4in_xing_in_r_mem_6_last; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_7_id = island_auto_axi4in_xing_in_r_mem_7_id; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_7_data = island_auto_axi4in_xing_in_r_mem_7_data; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_7_resp = island_auto_axi4in_xing_in_r_mem_7_resp; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_mem_7_last = island_auto_axi4in_xing_in_r_mem_7_last; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_widx = island_auto_axi4in_xing_in_r_widx; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_safe_widx_valid = island_auto_axi4in_xing_in_r_safe_widx_valid; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
  assign axi4asource_auto_out_r_safe_source_reset_n = island_auto_axi4in_xing_in_r_safe_source_reset_n; // @[LazyModule.scala 167:31:sifive.freedom.unleashed.DevKitU500FPGADesign_WithDevKit50MHz.fir@310819.4]
endmodule
