

module IBUFDS #(parameter   CAPACITANCE = "DONT_CARE",
                            DIFF_TERM = 0,
                            DQS_BIAS = 0,
                            IBUF_DELAY_VALUE = 0,
                            IBUF_LOW_PWR = 1,
                            IFD_DELAY_VALUE = "AUTO",
                            IOSTANDARD = "DEFAULT")(
   input I,
   input IB,
   output O
);


endmodule